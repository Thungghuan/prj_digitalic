module multiplier();

endmodule