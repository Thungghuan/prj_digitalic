module sin(sin_in, sin_out, sign);

input [9:0] sin_in;
output reg [12:0] sin_out;
output reg sign;

wire [1:0] high;
wire [7:0] low;

assign { high, low } = sin_in;

always @(*) begin
    case (high)
        2'b00: begin
            sign <= 1'b0;
            case (low)
                8'd000: sin_out <= 13'b0000000000000;
                8'd001: sin_out <= 13'b0000000011001;
                8'd002: sin_out <= 13'b0000000110010;
                8'd003: sin_out <= 13'b0000001001011;
                8'd004: sin_out <= 13'b0000001100101;
                8'd005: sin_out <= 13'b0000001111110;
                8'd006: sin_out <= 13'b0000010010111;
                8'd007: sin_out <= 13'b0000010110000;
                8'd008: sin_out <= 13'b0000011001001;
                8'd009: sin_out <= 13'b0000011100010;
                8'd010: sin_out <= 13'b0000011111011;
                8'd011: sin_out <= 13'b0000100010100;
                8'd012: sin_out <= 13'b0000100101101;
                8'd013: sin_out <= 13'b0000101000110;
                8'd014: sin_out <= 13'b0000101011111;
                8'd015: sin_out <= 13'b0000101111000;
                8'd016: sin_out <= 13'b0000110010001;
                8'd017: sin_out <= 13'b0000110101010;
                8'd018: sin_out <= 13'b0000111000011;
                8'd019: sin_out <= 13'b0000111011100;
                8'd020: sin_out <= 13'b0000111110101;
                8'd021: sin_out <= 13'b0001000001110;
                8'd022: sin_out <= 13'b0001000100111;
                8'd023: sin_out <= 13'b0001001000000;
                8'd024: sin_out <= 13'b0001001011001;
                8'd025: sin_out <= 13'b0001001110010;
                8'd026: sin_out <= 13'b0001010001011;
                8'd027: sin_out <= 13'b0001010100011;
                8'd028: sin_out <= 13'b0001010111100;
                8'd029: sin_out <= 13'b0001011010101;
                8'd030: sin_out <= 13'b0001011101110;
                8'd031: sin_out <= 13'b0001100000110;
                8'd032: sin_out <= 13'b0001100011111;
                8'd033: sin_out <= 13'b0001100111000;
                8'd034: sin_out <= 13'b0001101010000;
                8'd035: sin_out <= 13'b0001101101001;
                8'd036: sin_out <= 13'b0001110000001;
                8'd037: sin_out <= 13'b0001110011010;
                8'd038: sin_out <= 13'b0001110110010;
                8'd039: sin_out <= 13'b0001111001011;
                8'd040: sin_out <= 13'b0001111100011;
                8'd041: sin_out <= 13'b0001111111100;
                8'd042: sin_out <= 13'b0010000010100;
                8'd043: sin_out <= 13'b0010000101100;
                8'd044: sin_out <= 13'b0010001000100;
                8'd045: sin_out <= 13'b0010001011101;
                8'd046: sin_out <= 13'b0010001110101;
                8'd047: sin_out <= 13'b0010010001101;
                8'd048: sin_out <= 13'b0010010100101;
                8'd049: sin_out <= 13'b0010010111101;
                8'd050: sin_out <= 13'b0010011010101;
                8'd051: sin_out <= 13'b0010011101101;
                8'd052: sin_out <= 13'b0010100000101;
                8'd053: sin_out <= 13'b0010100011101;
                8'd054: sin_out <= 13'b0010100110100;
                8'd055: sin_out <= 13'b0010101001100;
                8'd056: sin_out <= 13'b0010101100100;
                8'd057: sin_out <= 13'b0010101111100;
                8'd058: sin_out <= 13'b0010110010011;
                8'd059: sin_out <= 13'b0010110101011;
                8'd060: sin_out <= 13'b0010111000010;
                8'd061: sin_out <= 13'b0010111011010;
                8'd062: sin_out <= 13'b0010111110001;
                8'd063: sin_out <= 13'b0011000001000;
                8'd064: sin_out <= 13'b0011000011111;
                8'd065: sin_out <= 13'b0011000110111;
                8'd066: sin_out <= 13'b0011001001110;
                8'd067: sin_out <= 13'b0011001100101;
                8'd068: sin_out <= 13'b0011001111100;
                8'd069: sin_out <= 13'b0011010010011;
                8'd070: sin_out <= 13'b0011010101010;
                8'd071: sin_out <= 13'b0011011000001;
                8'd072: sin_out <= 13'b0011011010111;
                8'd073: sin_out <= 13'b0011011101110;
                8'd074: sin_out <= 13'b0011100000101;
                8'd075: sin_out <= 13'b0011100011011;
                8'd076: sin_out <= 13'b0011100110010;
                8'd077: sin_out <= 13'b0011101001000;
                8'd078: sin_out <= 13'b0011101011110;
                8'd079: sin_out <= 13'b0011101110101;
                8'd080: sin_out <= 13'b0011110001011;
                8'd081: sin_out <= 13'b0011110100001;
                8'd082: sin_out <= 13'b0011110110111;
                8'd083: sin_out <= 13'b0011111001101;
                8'd084: sin_out <= 13'b0011111100011;
                8'd085: sin_out <= 13'b0011111111001;
                8'd086: sin_out <= 13'b0100000001110;
                8'd087: sin_out <= 13'b0100000100100;
                8'd088: sin_out <= 13'b0100000111010;
                8'd089: sin_out <= 13'b0100001001111;
                8'd090: sin_out <= 13'b0100001100101;
                8'd091: sin_out <= 13'b0100001111010;
                8'd092: sin_out <= 13'b0100010001111;
                8'd093: sin_out <= 13'b0100010100101;
                8'd094: sin_out <= 13'b0100010111010;
                8'd095: sin_out <= 13'b0100011001111;
                8'd096: sin_out <= 13'b0100011100100;
                8'd097: sin_out <= 13'b0100011111000;
                8'd098: sin_out <= 13'b0100100001101;
                8'd099: sin_out <= 13'b0100100100010;
                8'd100: sin_out <= 13'b0100100110111;
                8'd101: sin_out <= 13'b0100101001011;
                8'd102: sin_out <= 13'b0100101011111;
                8'd103: sin_out <= 13'b0100101110100;
                8'd104: sin_out <= 13'b0100110001000;
                8'd105: sin_out <= 13'b0100110011100;
                8'd106: sin_out <= 13'b0100110110000;
                8'd107: sin_out <= 13'b0100111000100;
                8'd108: sin_out <= 13'b0100111011000;
                8'd109: sin_out <= 13'b0100111101100;
                8'd110: sin_out <= 13'b0100111111111;
                8'd111: sin_out <= 13'b0101000010011;
                8'd112: sin_out <= 13'b0101000100110;
                8'd113: sin_out <= 13'b0101000111010;
                8'd114: sin_out <= 13'b0101001001101;
                8'd115: sin_out <= 13'b0101001100000;
                8'd116: sin_out <= 13'b0101001110011;
                8'd117: sin_out <= 13'b0101010000110;
                8'd118: sin_out <= 13'b0101010011001;
                8'd119: sin_out <= 13'b0101010101100;
                8'd120: sin_out <= 13'b0101010111111;
                8'd121: sin_out <= 13'b0101011010001;
                8'd122: sin_out <= 13'b0101011100100;
                8'd123: sin_out <= 13'b0101011110110;
                8'd124: sin_out <= 13'b0101100001000;
                8'd125: sin_out <= 13'b0101100011011;
                8'd126: sin_out <= 13'b0101100101101;
                8'd127: sin_out <= 13'b0101100111110;
                8'd128: sin_out <= 13'b0101101010000;
                8'd129: sin_out <= 13'b0101101100010;
                8'd130: sin_out <= 13'b0101101110100;
                8'd131: sin_out <= 13'b0101110000101;
                8'd132: sin_out <= 13'b0101110010111;
                8'd133: sin_out <= 13'b0101110101000;
                8'd134: sin_out <= 13'b0101110111001;
                8'd135: sin_out <= 13'b0101111001010;
                8'd136: sin_out <= 13'b0101111011011;
                8'd137: sin_out <= 13'b0101111101100;
                8'd138: sin_out <= 13'b0101111111100;
                8'd139: sin_out <= 13'b0110000001101;
                8'd140: sin_out <= 13'b0110000011110;
                8'd141: sin_out <= 13'b0110000101110;
                8'd142: sin_out <= 13'b0110000111110;
                8'd143: sin_out <= 13'b0110001001110;
                8'd144: sin_out <= 13'b0110001011110;
                8'd145: sin_out <= 13'b0110001101110;
                8'd146: sin_out <= 13'b0110001111110;
                8'd147: sin_out <= 13'b0110010001110;
                8'd148: sin_out <= 13'b0110010011101;
                8'd149: sin_out <= 13'b0110010101100;
                8'd150: sin_out <= 13'b0110010111100;
                8'd151: sin_out <= 13'b0110011001011;
                8'd152: sin_out <= 13'b0110011011010;
                8'd153: sin_out <= 13'b0110011101001;
                8'd154: sin_out <= 13'b0110011111000;
                8'd155: sin_out <= 13'b0110100000110;
                8'd156: sin_out <= 13'b0110100010101;
                8'd157: sin_out <= 13'b0110100100011;
                8'd158: sin_out <= 13'b0110100110010;
                8'd159: sin_out <= 13'b0110101000000;
                8'd160: sin_out <= 13'b0110101001110;
                8'd161: sin_out <= 13'b0110101011100;
                8'd162: sin_out <= 13'b0110101101001;
                8'd163: sin_out <= 13'b0110101110111;
                8'd164: sin_out <= 13'b0110110000101;
                8'd165: sin_out <= 13'b0110110010010;
                8'd166: sin_out <= 13'b0110110011111;
                8'd167: sin_out <= 13'b0110110101100;
                8'd168: sin_out <= 13'b0110110111001;
                8'd169: sin_out <= 13'b0110111000110;
                8'd170: sin_out <= 13'b0110111010011;
                8'd171: sin_out <= 13'b0110111011111;
                8'd172: sin_out <= 13'b0110111101100;
                8'd173: sin_out <= 13'b0110111111000;
                8'd174: sin_out <= 13'b0111000000100;
                8'd175: sin_out <= 13'b0111000010000;
                8'd176: sin_out <= 13'b0111000011100;
                8'd177: sin_out <= 13'b0111000101000;
                8'd178: sin_out <= 13'b0111000110100;
                8'd179: sin_out <= 13'b0111000111111;
                8'd180: sin_out <= 13'b0111001001011;
                8'd181: sin_out <= 13'b0111001010110;
                8'd182: sin_out <= 13'b0111001100001;
                8'd183: sin_out <= 13'b0111001101100;
                8'd184: sin_out <= 13'b0111001110111;
                8'd185: sin_out <= 13'b0111010000001;
                8'd186: sin_out <= 13'b0111010001100;
                8'd187: sin_out <= 13'b0111010010110;
                8'd188: sin_out <= 13'b0111010100001;
                8'd189: sin_out <= 13'b0111010101011;
                8'd190: sin_out <= 13'b0111010110101;
                8'd191: sin_out <= 13'b0111010111111;
                8'd192: sin_out <= 13'b0111011001000;
                8'd193: sin_out <= 13'b0111011010010;
                8'd194: sin_out <= 13'b0111011011011;
                8'd195: sin_out <= 13'b0111011100100;
                8'd196: sin_out <= 13'b0111011101110;
                8'd197: sin_out <= 13'b0111011110111;
                8'd198: sin_out <= 13'b0111011111111;
                8'd199: sin_out <= 13'b0111100001000;
                8'd200: sin_out <= 13'b0111100010001;
                8'd201: sin_out <= 13'b0111100011001;
                8'd202: sin_out <= 13'b0111100100001;
                8'd203: sin_out <= 13'b0111100101001;
                8'd204: sin_out <= 13'b0111100110001;
                8'd205: sin_out <= 13'b0111100111001;
                8'd206: sin_out <= 13'b0111101000001;
                8'd207: sin_out <= 13'b0111101001000;
                8'd208: sin_out <= 13'b0111101010000;
                8'd209: sin_out <= 13'b0111101010111;
                8'd210: sin_out <= 13'b0111101011110;
                8'd211: sin_out <= 13'b0111101100101;
                8'd212: sin_out <= 13'b0111101101100;
                8'd213: sin_out <= 13'b0111101110010;
                8'd214: sin_out <= 13'b0111101111001;
                8'd215: sin_out <= 13'b0111101111111;
                8'd216: sin_out <= 13'b0111110000101;
                8'd217: sin_out <= 13'b0111110001011;
                8'd218: sin_out <= 13'b0111110010001;
                8'd219: sin_out <= 13'b0111110010111;
                8'd220: sin_out <= 13'b0111110011100;
                8'd221: sin_out <= 13'b0111110100010;
                8'd222: sin_out <= 13'b0111110100111;
                8'd223: sin_out <= 13'b0111110101100;
                8'd224: sin_out <= 13'b0111110110001;
                8'd225: sin_out <= 13'b0111110110110;
                8'd226: sin_out <= 13'b0111110111011;
                8'd227: sin_out <= 13'b0111110111111;
                8'd228: sin_out <= 13'b0111111000100;
                8'd229: sin_out <= 13'b0111111001000;
                8'd230: sin_out <= 13'b0111111001100;
                8'd231: sin_out <= 13'b0111111010000;
                8'd232: sin_out <= 13'b0111111010100;
                8'd233: sin_out <= 13'b0111111010111;
                8'd234: sin_out <= 13'b0111111011011;
                8'd235: sin_out <= 13'b0111111011110;
                8'd236: sin_out <= 13'b0111111100001;
                8'd237: sin_out <= 13'b0111111100100;
                8'd238: sin_out <= 13'b0111111100111;
                8'd239: sin_out <= 13'b0111111101010;
                8'd240: sin_out <= 13'b0111111101100;
                8'd241: sin_out <= 13'b0111111101111;
                8'd242: sin_out <= 13'b0111111110001;
                8'd243: sin_out <= 13'b0111111110011;
                8'd244: sin_out <= 13'b0111111110101;
                8'd245: sin_out <= 13'b0111111110111;
                8'd246: sin_out <= 13'b0111111111000;
                8'd247: sin_out <= 13'b0111111111010;
                8'd248: sin_out <= 13'b0111111111011;
                8'd249: sin_out <= 13'b0111111111100;
                8'd250: sin_out <= 13'b0111111111101;
                8'd251: sin_out <= 13'b0111111111110;
                8'd252: sin_out <= 13'b0111111111111;
                8'd253: sin_out <= 13'b0111111111111;
                8'd254: sin_out <= 13'b1000000000000;
                8'd255: sin_out <= 13'b1000000000000;
            endcase
        end
        2'b01: begin
            sign <= 1'b0;
            case (low)
                8'd000: sin_out <= 13'b1000000000000;
                8'd001: sin_out <= 13'b1000000000000;
                8'd002: sin_out <= 13'b1000000000000;
                8'd003: sin_out <= 13'b0111111111111;
                8'd004: sin_out <= 13'b0111111111111;
                8'd005: sin_out <= 13'b0111111111110;
                8'd006: sin_out <= 13'b0111111111101;
                8'd007: sin_out <= 13'b0111111111100;
                8'd008: sin_out <= 13'b0111111111011;
                8'd009: sin_out <= 13'b0111111111010;
                8'd010: sin_out <= 13'b0111111111000;
                8'd011: sin_out <= 13'b0111111110111;
                8'd012: sin_out <= 13'b0111111110101;
                8'd013: sin_out <= 13'b0111111110011;
                8'd014: sin_out <= 13'b0111111110001;
                8'd015: sin_out <= 13'b0111111101111;
                8'd016: sin_out <= 13'b0111111101100;
                8'd017: sin_out <= 13'b0111111101010;
                8'd018: sin_out <= 13'b0111111100111;
                8'd019: sin_out <= 13'b0111111100100;
                8'd020: sin_out <= 13'b0111111100001;
                8'd021: sin_out <= 13'b0111111011110;
                8'd022: sin_out <= 13'b0111111011011;
                8'd023: sin_out <= 13'b0111111010111;
                8'd024: sin_out <= 13'b0111111010100;
                8'd025: sin_out <= 13'b0111111010000;
                8'd026: sin_out <= 13'b0111111001100;
                8'd027: sin_out <= 13'b0111111001000;
                8'd028: sin_out <= 13'b0111111000100;
                8'd029: sin_out <= 13'b0111110111111;
                8'd030: sin_out <= 13'b0111110111011;
                8'd031: sin_out <= 13'b0111110110110;
                8'd032: sin_out <= 13'b0111110110001;
                8'd033: sin_out <= 13'b0111110101100;
                8'd034: sin_out <= 13'b0111110100111;
                8'd035: sin_out <= 13'b0111110100010;
                8'd036: sin_out <= 13'b0111110011100;
                8'd037: sin_out <= 13'b0111110010111;
                8'd038: sin_out <= 13'b0111110010001;
                8'd039: sin_out <= 13'b0111110001011;
                8'd040: sin_out <= 13'b0111110000101;
                8'd041: sin_out <= 13'b0111101111111;
                8'd042: sin_out <= 13'b0111101111001;
                8'd043: sin_out <= 13'b0111101110010;
                8'd044: sin_out <= 13'b0111101101100;
                8'd045: sin_out <= 13'b0111101100101;
                8'd046: sin_out <= 13'b0111101011110;
                8'd047: sin_out <= 13'b0111101010111;
                8'd048: sin_out <= 13'b0111101010000;
                8'd049: sin_out <= 13'b0111101001000;
                8'd050: sin_out <= 13'b0111101000001;
                8'd051: sin_out <= 13'b0111100111001;
                8'd052: sin_out <= 13'b0111100110001;
                8'd053: sin_out <= 13'b0111100101001;
                8'd054: sin_out <= 13'b0111100100001;
                8'd055: sin_out <= 13'b0111100011001;
                8'd056: sin_out <= 13'b0111100010001;
                8'd057: sin_out <= 13'b0111100001000;
                8'd058: sin_out <= 13'b0111011111111;
                8'd059: sin_out <= 13'b0111011110111;
                8'd060: sin_out <= 13'b0111011101110;
                8'd061: sin_out <= 13'b0111011100100;
                8'd062: sin_out <= 13'b0111011011011;
                8'd063: sin_out <= 13'b0111011010010;
                8'd064: sin_out <= 13'b0111011001000;
                8'd065: sin_out <= 13'b0111010111111;
                8'd066: sin_out <= 13'b0111010110101;
                8'd067: sin_out <= 13'b0111010101011;
                8'd068: sin_out <= 13'b0111010100001;
                8'd069: sin_out <= 13'b0111010010110;
                8'd070: sin_out <= 13'b0111010001100;
                8'd071: sin_out <= 13'b0111010000001;
                8'd072: sin_out <= 13'b0111001110111;
                8'd073: sin_out <= 13'b0111001101100;
                8'd074: sin_out <= 13'b0111001100001;
                8'd075: sin_out <= 13'b0111001010110;
                8'd076: sin_out <= 13'b0111001001011;
                8'd077: sin_out <= 13'b0111000111111;
                8'd078: sin_out <= 13'b0111000110100;
                8'd079: sin_out <= 13'b0111000101000;
                8'd080: sin_out <= 13'b0111000011100;
                8'd081: sin_out <= 13'b0111000010000;
                8'd082: sin_out <= 13'b0111000000100;
                8'd083: sin_out <= 13'b0110111111000;
                8'd084: sin_out <= 13'b0110111101100;
                8'd085: sin_out <= 13'b0110111011111;
                8'd086: sin_out <= 13'b0110111010011;
                8'd087: sin_out <= 13'b0110111000110;
                8'd088: sin_out <= 13'b0110110111001;
                8'd089: sin_out <= 13'b0110110101100;
                8'd090: sin_out <= 13'b0110110011111;
                8'd091: sin_out <= 13'b0110110010010;
                8'd092: sin_out <= 13'b0110110000101;
                8'd093: sin_out <= 13'b0110101110111;
                8'd094: sin_out <= 13'b0110101101001;
                8'd095: sin_out <= 13'b0110101011100;
                8'd096: sin_out <= 13'b0110101001110;
                8'd097: sin_out <= 13'b0110101000000;
                8'd098: sin_out <= 13'b0110100110010;
                8'd099: sin_out <= 13'b0110100100011;
                8'd100: sin_out <= 13'b0110100010101;
                8'd101: sin_out <= 13'b0110100000110;
                8'd102: sin_out <= 13'b0110011111000;
                8'd103: sin_out <= 13'b0110011101001;
                8'd104: sin_out <= 13'b0110011011010;
                8'd105: sin_out <= 13'b0110011001011;
                8'd106: sin_out <= 13'b0110010111100;
                8'd107: sin_out <= 13'b0110010101100;
                8'd108: sin_out <= 13'b0110010011101;
                8'd109: sin_out <= 13'b0110010001110;
                8'd110: sin_out <= 13'b0110001111110;
                8'd111: sin_out <= 13'b0110001101110;
                8'd112: sin_out <= 13'b0110001011110;
                8'd113: sin_out <= 13'b0110001001110;
                8'd114: sin_out <= 13'b0110000111110;
                8'd115: sin_out <= 13'b0110000101110;
                8'd116: sin_out <= 13'b0110000011110;
                8'd117: sin_out <= 13'b0110000001101;
                8'd118: sin_out <= 13'b0101111111100;
                8'd119: sin_out <= 13'b0101111101100;
                8'd120: sin_out <= 13'b0101111011011;
                8'd121: sin_out <= 13'b0101111001010;
                8'd122: sin_out <= 13'b0101110111001;
                8'd123: sin_out <= 13'b0101110101000;
                8'd124: sin_out <= 13'b0101110010111;
                8'd125: sin_out <= 13'b0101110000101;
                8'd126: sin_out <= 13'b0101101110100;
                8'd127: sin_out <= 13'b0101101100010;
                8'd128: sin_out <= 13'b0101101010000;
                8'd129: sin_out <= 13'b0101100111110;
                8'd130: sin_out <= 13'b0101100101101;
                8'd131: sin_out <= 13'b0101100011011;
                8'd132: sin_out <= 13'b0101100001000;
                8'd133: sin_out <= 13'b0101011110110;
                8'd134: sin_out <= 13'b0101011100100;
                8'd135: sin_out <= 13'b0101011010001;
                8'd136: sin_out <= 13'b0101010111111;
                8'd137: sin_out <= 13'b0101010101100;
                8'd138: sin_out <= 13'b0101010011001;
                8'd139: sin_out <= 13'b0101010000110;
                8'd140: sin_out <= 13'b0101001110011;
                8'd141: sin_out <= 13'b0101001100000;
                8'd142: sin_out <= 13'b0101001001101;
                8'd143: sin_out <= 13'b0101000111010;
                8'd144: sin_out <= 13'b0101000100110;
                8'd145: sin_out <= 13'b0101000010011;
                8'd146: sin_out <= 13'b0100111111111;
                8'd147: sin_out <= 13'b0100111101100;
                8'd148: sin_out <= 13'b0100111011000;
                8'd149: sin_out <= 13'b0100111000100;
                8'd150: sin_out <= 13'b0100110110000;
                8'd151: sin_out <= 13'b0100110011100;
                8'd152: sin_out <= 13'b0100110001000;
                8'd153: sin_out <= 13'b0100101110100;
                8'd154: sin_out <= 13'b0100101011111;
                8'd155: sin_out <= 13'b0100101001011;
                8'd156: sin_out <= 13'b0100100110111;
                8'd157: sin_out <= 13'b0100100100010;
                8'd158: sin_out <= 13'b0100100001101;
                8'd159: sin_out <= 13'b0100011111000;
                8'd160: sin_out <= 13'b0100011100100;
                8'd161: sin_out <= 13'b0100011001111;
                8'd162: sin_out <= 13'b0100010111010;
                8'd163: sin_out <= 13'b0100010100101;
                8'd164: sin_out <= 13'b0100010001111;
                8'd165: sin_out <= 13'b0100001111010;
                8'd166: sin_out <= 13'b0100001100101;
                8'd167: sin_out <= 13'b0100001001111;
                8'd168: sin_out <= 13'b0100000111010;
                8'd169: sin_out <= 13'b0100000100100;
                8'd170: sin_out <= 13'b0100000001110;
                8'd171: sin_out <= 13'b0011111111001;
                8'd172: sin_out <= 13'b0011111100011;
                8'd173: sin_out <= 13'b0011111001101;
                8'd174: sin_out <= 13'b0011110110111;
                8'd175: sin_out <= 13'b0011110100001;
                8'd176: sin_out <= 13'b0011110001011;
                8'd177: sin_out <= 13'b0011101110101;
                8'd178: sin_out <= 13'b0011101011110;
                8'd179: sin_out <= 13'b0011101001000;
                8'd180: sin_out <= 13'b0011100110010;
                8'd181: sin_out <= 13'b0011100011011;
                8'd182: sin_out <= 13'b0011100000101;
                8'd183: sin_out <= 13'b0011011101110;
                8'd184: sin_out <= 13'b0011011010111;
                8'd185: sin_out <= 13'b0011011000001;
                8'd186: sin_out <= 13'b0011010101010;
                8'd187: sin_out <= 13'b0011010010011;
                8'd188: sin_out <= 13'b0011001111100;
                8'd189: sin_out <= 13'b0011001100101;
                8'd190: sin_out <= 13'b0011001001110;
                8'd191: sin_out <= 13'b0011000110111;
                8'd192: sin_out <= 13'b0011000011111;
                8'd193: sin_out <= 13'b0011000001000;
                8'd194: sin_out <= 13'b0010111110001;
                8'd195: sin_out <= 13'b0010111011010;
                8'd196: sin_out <= 13'b0010111000010;
                8'd197: sin_out <= 13'b0010110101011;
                8'd198: sin_out <= 13'b0010110010011;
                8'd199: sin_out <= 13'b0010101111100;
                8'd200: sin_out <= 13'b0010101100100;
                8'd201: sin_out <= 13'b0010101001100;
                8'd202: sin_out <= 13'b0010100110100;
                8'd203: sin_out <= 13'b0010100011101;
                8'd204: sin_out <= 13'b0010100000101;
                8'd205: sin_out <= 13'b0010011101101;
                8'd206: sin_out <= 13'b0010011010101;
                8'd207: sin_out <= 13'b0010010111101;
                8'd208: sin_out <= 13'b0010010100101;
                8'd209: sin_out <= 13'b0010010001101;
                8'd210: sin_out <= 13'b0010001110101;
                8'd211: sin_out <= 13'b0010001011101;
                8'd212: sin_out <= 13'b0010001000100;
                8'd213: sin_out <= 13'b0010000101100;
                8'd214: sin_out <= 13'b0010000010100;
                8'd215: sin_out <= 13'b0001111111100;
                8'd216: sin_out <= 13'b0001111100011;
                8'd217: sin_out <= 13'b0001111001011;
                8'd218: sin_out <= 13'b0001110110010;
                8'd219: sin_out <= 13'b0001110011010;
                8'd220: sin_out <= 13'b0001110000001;
                8'd221: sin_out <= 13'b0001101101001;
                8'd222: sin_out <= 13'b0001101010000;
                8'd223: sin_out <= 13'b0001100111000;
                8'd224: sin_out <= 13'b0001100011111;
                8'd225: sin_out <= 13'b0001100000110;
                8'd226: sin_out <= 13'b0001011101110;
                8'd227: sin_out <= 13'b0001011010101;
                8'd228: sin_out <= 13'b0001010111100;
                8'd229: sin_out <= 13'b0001010100011;
                8'd230: sin_out <= 13'b0001010001011;
                8'd231: sin_out <= 13'b0001001110010;
                8'd232: sin_out <= 13'b0001001011001;
                8'd233: sin_out <= 13'b0001001000000;
                8'd234: sin_out <= 13'b0001000100111;
                8'd235: sin_out <= 13'b0001000001110;
                8'd236: sin_out <= 13'b0000111110101;
                8'd237: sin_out <= 13'b0000111011100;
                8'd238: sin_out <= 13'b0000111000011;
                8'd239: sin_out <= 13'b0000110101010;
                8'd240: sin_out <= 13'b0000110010001;
                8'd241: sin_out <= 13'b0000101111000;
                8'd242: sin_out <= 13'b0000101011111;
                8'd243: sin_out <= 13'b0000101000110;
                8'd244: sin_out <= 13'b0000100101101;
                8'd245: sin_out <= 13'b0000100010100;
                8'd246: sin_out <= 13'b0000011111011;
                8'd247: sin_out <= 13'b0000011100010;
                8'd248: sin_out <= 13'b0000011001001;
                8'd249: sin_out <= 13'b0000010110000;
                8'd250: sin_out <= 13'b0000010010111;
                8'd251: sin_out <= 13'b0000001111110;
                8'd252: sin_out <= 13'b0000001100101;
                8'd253: sin_out <= 13'b0000001001011;
                8'd254: sin_out <= 13'b0000000110010;
                8'd255: sin_out <= 13'b0000000011001;
            endcase
        end
        2'b10: begin
            sign <= 1'b1;
            case (low)
                8'd000: sin_out <= 13'b0000000000000;
                8'd001: sin_out <= 13'b0000000011001;
                8'd002: sin_out <= 13'b0000000110010;
                8'd003: sin_out <= 13'b0000001001011;
                8'd004: sin_out <= 13'b0000001100101;
                8'd005: sin_out <= 13'b0000001111110;
                8'd006: sin_out <= 13'b0000010010111;
                8'd007: sin_out <= 13'b0000010110000;
                8'd008: sin_out <= 13'b0000011001001;
                8'd009: sin_out <= 13'b0000011100010;
                8'd010: sin_out <= 13'b0000011111011;
                8'd011: sin_out <= 13'b0000100010100;
                8'd012: sin_out <= 13'b0000100101101;
                8'd013: sin_out <= 13'b0000101000110;
                8'd014: sin_out <= 13'b0000101011111;
                8'd015: sin_out <= 13'b0000101111000;
                8'd016: sin_out <= 13'b0000110010001;
                8'd017: sin_out <= 13'b0000110101010;
                8'd018: sin_out <= 13'b0000111000011;
                8'd019: sin_out <= 13'b0000111011100;
                8'd020: sin_out <= 13'b0000111110101;
                8'd021: sin_out <= 13'b0001000001110;
                8'd022: sin_out <= 13'b0001000100111;
                8'd023: sin_out <= 13'b0001001000000;
                8'd024: sin_out <= 13'b0001001011001;
                8'd025: sin_out <= 13'b0001001110010;
                8'd026: sin_out <= 13'b0001010001011;
                8'd027: sin_out <= 13'b0001010100011;
                8'd028: sin_out <= 13'b0001010111100;
                8'd029: sin_out <= 13'b0001011010101;
                8'd030: sin_out <= 13'b0001011101110;
                8'd031: sin_out <= 13'b0001100000110;
                8'd032: sin_out <= 13'b0001100011111;
                8'd033: sin_out <= 13'b0001100111000;
                8'd034: sin_out <= 13'b0001101010000;
                8'd035: sin_out <= 13'b0001101101001;
                8'd036: sin_out <= 13'b0001110000001;
                8'd037: sin_out <= 13'b0001110011010;
                8'd038: sin_out <= 13'b0001110110010;
                8'd039: sin_out <= 13'b0001111001011;
                8'd040: sin_out <= 13'b0001111100011;
                8'd041: sin_out <= 13'b0001111111100;
                8'd042: sin_out <= 13'b0010000010100;
                8'd043: sin_out <= 13'b0010000101100;
                8'd044: sin_out <= 13'b0010001000100;
                8'd045: sin_out <= 13'b0010001011101;
                8'd046: sin_out <= 13'b0010001110101;
                8'd047: sin_out <= 13'b0010010001101;
                8'd048: sin_out <= 13'b0010010100101;
                8'd049: sin_out <= 13'b0010010111101;
                8'd050: sin_out <= 13'b0010011010101;
                8'd051: sin_out <= 13'b0010011101101;
                8'd052: sin_out <= 13'b0010100000101;
                8'd053: sin_out <= 13'b0010100011101;
                8'd054: sin_out <= 13'b0010100110100;
                8'd055: sin_out <= 13'b0010101001100;
                8'd056: sin_out <= 13'b0010101100100;
                8'd057: sin_out <= 13'b0010101111100;
                8'd058: sin_out <= 13'b0010110010011;
                8'd059: sin_out <= 13'b0010110101011;
                8'd060: sin_out <= 13'b0010111000010;
                8'd061: sin_out <= 13'b0010111011010;
                8'd062: sin_out <= 13'b0010111110001;
                8'd063: sin_out <= 13'b0011000001000;
                8'd064: sin_out <= 13'b0011000011111;
                8'd065: sin_out <= 13'b0011000110111;
                8'd066: sin_out <= 13'b0011001001110;
                8'd067: sin_out <= 13'b0011001100101;
                8'd068: sin_out <= 13'b0011001111100;
                8'd069: sin_out <= 13'b0011010010011;
                8'd070: sin_out <= 13'b0011010101010;
                8'd071: sin_out <= 13'b0011011000001;
                8'd072: sin_out <= 13'b0011011010111;
                8'd073: sin_out <= 13'b0011011101110;
                8'd074: sin_out <= 13'b0011100000101;
                8'd075: sin_out <= 13'b0011100011011;
                8'd076: sin_out <= 13'b0011100110010;
                8'd077: sin_out <= 13'b0011101001000;
                8'd078: sin_out <= 13'b0011101011110;
                8'd079: sin_out <= 13'b0011101110101;
                8'd080: sin_out <= 13'b0011110001011;
                8'd081: sin_out <= 13'b0011110100001;
                8'd082: sin_out <= 13'b0011110110111;
                8'd083: sin_out <= 13'b0011111001101;
                8'd084: sin_out <= 13'b0011111100011;
                8'd085: sin_out <= 13'b0011111111001;
                8'd086: sin_out <= 13'b0100000001110;
                8'd087: sin_out <= 13'b0100000100100;
                8'd088: sin_out <= 13'b0100000111010;
                8'd089: sin_out <= 13'b0100001001111;
                8'd090: sin_out <= 13'b0100001100101;
                8'd091: sin_out <= 13'b0100001111010;
                8'd092: sin_out <= 13'b0100010001111;
                8'd093: sin_out <= 13'b0100010100101;
                8'd094: sin_out <= 13'b0100010111010;
                8'd095: sin_out <= 13'b0100011001111;
                8'd096: sin_out <= 13'b0100011100100;
                8'd097: sin_out <= 13'b0100011111000;
                8'd098: sin_out <= 13'b0100100001101;
                8'd099: sin_out <= 13'b0100100100010;
                8'd100: sin_out <= 13'b0100100110111;
                8'd101: sin_out <= 13'b0100101001011;
                8'd102: sin_out <= 13'b0100101011111;
                8'd103: sin_out <= 13'b0100101110100;
                8'd104: sin_out <= 13'b0100110001000;
                8'd105: sin_out <= 13'b0100110011100;
                8'd106: sin_out <= 13'b0100110110000;
                8'd107: sin_out <= 13'b0100111000100;
                8'd108: sin_out <= 13'b0100111011000;
                8'd109: sin_out <= 13'b0100111101100;
                8'd110: sin_out <= 13'b0100111111111;
                8'd111: sin_out <= 13'b0101000010011;
                8'd112: sin_out <= 13'b0101000100110;
                8'd113: sin_out <= 13'b0101000111010;
                8'd114: sin_out <= 13'b0101001001101;
                8'd115: sin_out <= 13'b0101001100000;
                8'd116: sin_out <= 13'b0101001110011;
                8'd117: sin_out <= 13'b0101010000110;
                8'd118: sin_out <= 13'b0101010011001;
                8'd119: sin_out <= 13'b0101010101100;
                8'd120: sin_out <= 13'b0101010111111;
                8'd121: sin_out <= 13'b0101011010001;
                8'd122: sin_out <= 13'b0101011100100;
                8'd123: sin_out <= 13'b0101011110110;
                8'd124: sin_out <= 13'b0101100001000;
                8'd125: sin_out <= 13'b0101100011011;
                8'd126: sin_out <= 13'b0101100101101;
                8'd127: sin_out <= 13'b0101100111110;
                8'd128: sin_out <= 13'b0101101010000;
                8'd129: sin_out <= 13'b0101101100010;
                8'd130: sin_out <= 13'b0101101110100;
                8'd131: sin_out <= 13'b0101110000101;
                8'd132: sin_out <= 13'b0101110010111;
                8'd133: sin_out <= 13'b0101110101000;
                8'd134: sin_out <= 13'b0101110111001;
                8'd135: sin_out <= 13'b0101111001010;
                8'd136: sin_out <= 13'b0101111011011;
                8'd137: sin_out <= 13'b0101111101100;
                8'd138: sin_out <= 13'b0101111111100;
                8'd139: sin_out <= 13'b0110000001101;
                8'd140: sin_out <= 13'b0110000011110;
                8'd141: sin_out <= 13'b0110000101110;
                8'd142: sin_out <= 13'b0110000111110;
                8'd143: sin_out <= 13'b0110001001110;
                8'd144: sin_out <= 13'b0110001011110;
                8'd145: sin_out <= 13'b0110001101110;
                8'd146: sin_out <= 13'b0110001111110;
                8'd147: sin_out <= 13'b0110010001110;
                8'd148: sin_out <= 13'b0110010011101;
                8'd149: sin_out <= 13'b0110010101100;
                8'd150: sin_out <= 13'b0110010111100;
                8'd151: sin_out <= 13'b0110011001011;
                8'd152: sin_out <= 13'b0110011011010;
                8'd153: sin_out <= 13'b0110011101001;
                8'd154: sin_out <= 13'b0110011111000;
                8'd155: sin_out <= 13'b0110100000110;
                8'd156: sin_out <= 13'b0110100010101;
                8'd157: sin_out <= 13'b0110100100011;
                8'd158: sin_out <= 13'b0110100110010;
                8'd159: sin_out <= 13'b0110101000000;
                8'd160: sin_out <= 13'b0110101001110;
                8'd161: sin_out <= 13'b0110101011100;
                8'd162: sin_out <= 13'b0110101101001;
                8'd163: sin_out <= 13'b0110101110111;
                8'd164: sin_out <= 13'b0110110000101;
                8'd165: sin_out <= 13'b0110110010010;
                8'd166: sin_out <= 13'b0110110011111;
                8'd167: sin_out <= 13'b0110110101100;
                8'd168: sin_out <= 13'b0110110111001;
                8'd169: sin_out <= 13'b0110111000110;
                8'd170: sin_out <= 13'b0110111010011;
                8'd171: sin_out <= 13'b0110111011111;
                8'd172: sin_out <= 13'b0110111101100;
                8'd173: sin_out <= 13'b0110111111000;
                8'd174: sin_out <= 13'b0111000000100;
                8'd175: sin_out <= 13'b0111000010000;
                8'd176: sin_out <= 13'b0111000011100;
                8'd177: sin_out <= 13'b0111000101000;
                8'd178: sin_out <= 13'b0111000110100;
                8'd179: sin_out <= 13'b0111000111111;
                8'd180: sin_out <= 13'b0111001001011;
                8'd181: sin_out <= 13'b0111001010110;
                8'd182: sin_out <= 13'b0111001100001;
                8'd183: sin_out <= 13'b0111001101100;
                8'd184: sin_out <= 13'b0111001110111;
                8'd185: sin_out <= 13'b0111010000001;
                8'd186: sin_out <= 13'b0111010001100;
                8'd187: sin_out <= 13'b0111010010110;
                8'd188: sin_out <= 13'b0111010100001;
                8'd189: sin_out <= 13'b0111010101011;
                8'd190: sin_out <= 13'b0111010110101;
                8'd191: sin_out <= 13'b0111010111111;
                8'd192: sin_out <= 13'b0111011001000;
                8'd193: sin_out <= 13'b0111011010010;
                8'd194: sin_out <= 13'b0111011011011;
                8'd195: sin_out <= 13'b0111011100100;
                8'd196: sin_out <= 13'b0111011101110;
                8'd197: sin_out <= 13'b0111011110111;
                8'd198: sin_out <= 13'b0111011111111;
                8'd199: sin_out <= 13'b0111100001000;
                8'd200: sin_out <= 13'b0111100010001;
                8'd201: sin_out <= 13'b0111100011001;
                8'd202: sin_out <= 13'b0111100100001;
                8'd203: sin_out <= 13'b0111100101001;
                8'd204: sin_out <= 13'b0111100110001;
                8'd205: sin_out <= 13'b0111100111001;
                8'd206: sin_out <= 13'b0111101000001;
                8'd207: sin_out <= 13'b0111101001000;
                8'd208: sin_out <= 13'b0111101010000;
                8'd209: sin_out <= 13'b0111101010111;
                8'd210: sin_out <= 13'b0111101011110;
                8'd211: sin_out <= 13'b0111101100101;
                8'd212: sin_out <= 13'b0111101101100;
                8'd213: sin_out <= 13'b0111101110010;
                8'd214: sin_out <= 13'b0111101111001;
                8'd215: sin_out <= 13'b0111101111111;
                8'd216: sin_out <= 13'b0111110000101;
                8'd217: sin_out <= 13'b0111110001011;
                8'd218: sin_out <= 13'b0111110010001;
                8'd219: sin_out <= 13'b0111110010111;
                8'd220: sin_out <= 13'b0111110011100;
                8'd221: sin_out <= 13'b0111110100010;
                8'd222: sin_out <= 13'b0111110100111;
                8'd223: sin_out <= 13'b0111110101100;
                8'd224: sin_out <= 13'b0111110110001;
                8'd225: sin_out <= 13'b0111110110110;
                8'd226: sin_out <= 13'b0111110111011;
                8'd227: sin_out <= 13'b0111110111111;
                8'd228: sin_out <= 13'b0111111000100;
                8'd229: sin_out <= 13'b0111111001000;
                8'd230: sin_out <= 13'b0111111001100;
                8'd231: sin_out <= 13'b0111111010000;
                8'd232: sin_out <= 13'b0111111010100;
                8'd233: sin_out <= 13'b0111111010111;
                8'd234: sin_out <= 13'b0111111011011;
                8'd235: sin_out <= 13'b0111111011110;
                8'd236: sin_out <= 13'b0111111100001;
                8'd237: sin_out <= 13'b0111111100100;
                8'd238: sin_out <= 13'b0111111100111;
                8'd239: sin_out <= 13'b0111111101010;
                8'd240: sin_out <= 13'b0111111101100;
                8'd241: sin_out <= 13'b0111111101111;
                8'd242: sin_out <= 13'b0111111110001;
                8'd243: sin_out <= 13'b0111111110011;
                8'd244: sin_out <= 13'b0111111110101;
                8'd245: sin_out <= 13'b0111111110111;
                8'd246: sin_out <= 13'b0111111111000;
                8'd247: sin_out <= 13'b0111111111010;
                8'd248: sin_out <= 13'b0111111111011;
                8'd249: sin_out <= 13'b0111111111100;
                8'd250: sin_out <= 13'b0111111111101;
                8'd251: sin_out <= 13'b0111111111110;
                8'd252: sin_out <= 13'b0111111111111;
                8'd253: sin_out <= 13'b0111111111111;
                8'd254: sin_out <= 13'b1000000000000;
                8'd255: sin_out <= 13'b1000000000000;
            endcase
        end
        2'b11: begin
            sign <= 1'b1;
            case (low)
                8'd000: sin_out <= 13'b1000000000000;
                8'd001: sin_out <= 13'b1000000000000;
                8'd002: sin_out <= 13'b1000000000000;
                8'd003: sin_out <= 13'b0111111111111;
                8'd004: sin_out <= 13'b0111111111111;
                8'd005: sin_out <= 13'b0111111111110;
                8'd006: sin_out <= 13'b0111111111101;
                8'd007: sin_out <= 13'b0111111111100;
                8'd008: sin_out <= 13'b0111111111011;
                8'd009: sin_out <= 13'b0111111111010;
                8'd010: sin_out <= 13'b0111111111000;
                8'd011: sin_out <= 13'b0111111110111;
                8'd012: sin_out <= 13'b0111111110101;
                8'd013: sin_out <= 13'b0111111110011;
                8'd014: sin_out <= 13'b0111111110001;
                8'd015: sin_out <= 13'b0111111101111;
                8'd016: sin_out <= 13'b0111111101100;
                8'd017: sin_out <= 13'b0111111101010;
                8'd018: sin_out <= 13'b0111111100111;
                8'd019: sin_out <= 13'b0111111100100;
                8'd020: sin_out <= 13'b0111111100001;
                8'd021: sin_out <= 13'b0111111011110;
                8'd022: sin_out <= 13'b0111111011011;
                8'd023: sin_out <= 13'b0111111010111;
                8'd024: sin_out <= 13'b0111111010100;
                8'd025: sin_out <= 13'b0111111010000;
                8'd026: sin_out <= 13'b0111111001100;
                8'd027: sin_out <= 13'b0111111001000;
                8'd028: sin_out <= 13'b0111111000100;
                8'd029: sin_out <= 13'b0111110111111;
                8'd030: sin_out <= 13'b0111110111011;
                8'd031: sin_out <= 13'b0111110110110;
                8'd032: sin_out <= 13'b0111110110001;
                8'd033: sin_out <= 13'b0111110101100;
                8'd034: sin_out <= 13'b0111110100111;
                8'd035: sin_out <= 13'b0111110100010;
                8'd036: sin_out <= 13'b0111110011100;
                8'd037: sin_out <= 13'b0111110010111;
                8'd038: sin_out <= 13'b0111110010001;
                8'd039: sin_out <= 13'b0111110001011;
                8'd040: sin_out <= 13'b0111110000101;
                8'd041: sin_out <= 13'b0111101111111;
                8'd042: sin_out <= 13'b0111101111001;
                8'd043: sin_out <= 13'b0111101110010;
                8'd044: sin_out <= 13'b0111101101100;
                8'd045: sin_out <= 13'b0111101100101;
                8'd046: sin_out <= 13'b0111101011110;
                8'd047: sin_out <= 13'b0111101010111;
                8'd048: sin_out <= 13'b0111101010000;
                8'd049: sin_out <= 13'b0111101001000;
                8'd050: sin_out <= 13'b0111101000001;
                8'd051: sin_out <= 13'b0111100111001;
                8'd052: sin_out <= 13'b0111100110001;
                8'd053: sin_out <= 13'b0111100101001;
                8'd054: sin_out <= 13'b0111100100001;
                8'd055: sin_out <= 13'b0111100011001;
                8'd056: sin_out <= 13'b0111100010001;
                8'd057: sin_out <= 13'b0111100001000;
                8'd058: sin_out <= 13'b0111011111111;
                8'd059: sin_out <= 13'b0111011110111;
                8'd060: sin_out <= 13'b0111011101110;
                8'd061: sin_out <= 13'b0111011100100;
                8'd062: sin_out <= 13'b0111011011011;
                8'd063: sin_out <= 13'b0111011010010;
                8'd064: sin_out <= 13'b0111011001000;
                8'd065: sin_out <= 13'b0111010111111;
                8'd066: sin_out <= 13'b0111010110101;
                8'd067: sin_out <= 13'b0111010101011;
                8'd068: sin_out <= 13'b0111010100001;
                8'd069: sin_out <= 13'b0111010010110;
                8'd070: sin_out <= 13'b0111010001100;
                8'd071: sin_out <= 13'b0111010000001;
                8'd072: sin_out <= 13'b0111001110111;
                8'd073: sin_out <= 13'b0111001101100;
                8'd074: sin_out <= 13'b0111001100001;
                8'd075: sin_out <= 13'b0111001010110;
                8'd076: sin_out <= 13'b0111001001011;
                8'd077: sin_out <= 13'b0111000111111;
                8'd078: sin_out <= 13'b0111000110100;
                8'd079: sin_out <= 13'b0111000101000;
                8'd080: sin_out <= 13'b0111000011100;
                8'd081: sin_out <= 13'b0111000010000;
                8'd082: sin_out <= 13'b0111000000100;
                8'd083: sin_out <= 13'b0110111111000;
                8'd084: sin_out <= 13'b0110111101100;
                8'd085: sin_out <= 13'b0110111011111;
                8'd086: sin_out <= 13'b0110111010011;
                8'd087: sin_out <= 13'b0110111000110;
                8'd088: sin_out <= 13'b0110110111001;
                8'd089: sin_out <= 13'b0110110101100;
                8'd090: sin_out <= 13'b0110110011111;
                8'd091: sin_out <= 13'b0110110010010;
                8'd092: sin_out <= 13'b0110110000101;
                8'd093: sin_out <= 13'b0110101110111;
                8'd094: sin_out <= 13'b0110101101001;
                8'd095: sin_out <= 13'b0110101011100;
                8'd096: sin_out <= 13'b0110101001110;
                8'd097: sin_out <= 13'b0110101000000;
                8'd098: sin_out <= 13'b0110100110010;
                8'd099: sin_out <= 13'b0110100100011;
                8'd100: sin_out <= 13'b0110100010101;
                8'd101: sin_out <= 13'b0110100000110;
                8'd102: sin_out <= 13'b0110011111000;
                8'd103: sin_out <= 13'b0110011101001;
                8'd104: sin_out <= 13'b0110011011010;
                8'd105: sin_out <= 13'b0110011001011;
                8'd106: sin_out <= 13'b0110010111100;
                8'd107: sin_out <= 13'b0110010101100;
                8'd108: sin_out <= 13'b0110010011101;
                8'd109: sin_out <= 13'b0110010001110;
                8'd110: sin_out <= 13'b0110001111110;
                8'd111: sin_out <= 13'b0110001101110;
                8'd112: sin_out <= 13'b0110001011110;
                8'd113: sin_out <= 13'b0110001001110;
                8'd114: sin_out <= 13'b0110000111110;
                8'd115: sin_out <= 13'b0110000101110;
                8'd116: sin_out <= 13'b0110000011110;
                8'd117: sin_out <= 13'b0110000001101;
                8'd118: sin_out <= 13'b0101111111100;
                8'd119: sin_out <= 13'b0101111101100;
                8'd120: sin_out <= 13'b0101111011011;
                8'd121: sin_out <= 13'b0101111001010;
                8'd122: sin_out <= 13'b0101110111001;
                8'd123: sin_out <= 13'b0101110101000;
                8'd124: sin_out <= 13'b0101110010111;
                8'd125: sin_out <= 13'b0101110000101;
                8'd126: sin_out <= 13'b0101101110100;
                8'd127: sin_out <= 13'b0101101100010;
                8'd128: sin_out <= 13'b0101101010000;
                8'd129: sin_out <= 13'b0101100111110;
                8'd130: sin_out <= 13'b0101100101101;
                8'd131: sin_out <= 13'b0101100011011;
                8'd132: sin_out <= 13'b0101100001000;
                8'd133: sin_out <= 13'b0101011110110;
                8'd134: sin_out <= 13'b0101011100100;
                8'd135: sin_out <= 13'b0101011010001;
                8'd136: sin_out <= 13'b0101010111111;
                8'd137: sin_out <= 13'b0101010101100;
                8'd138: sin_out <= 13'b0101010011001;
                8'd139: sin_out <= 13'b0101010000110;
                8'd140: sin_out <= 13'b0101001110011;
                8'd141: sin_out <= 13'b0101001100000;
                8'd142: sin_out <= 13'b0101001001101;
                8'd143: sin_out <= 13'b0101000111010;
                8'd144: sin_out <= 13'b0101000100110;
                8'd145: sin_out <= 13'b0101000010011;
                8'd146: sin_out <= 13'b0100111111111;
                8'd147: sin_out <= 13'b0100111101100;
                8'd148: sin_out <= 13'b0100111011000;
                8'd149: sin_out <= 13'b0100111000100;
                8'd150: sin_out <= 13'b0100110110000;
                8'd151: sin_out <= 13'b0100110011100;
                8'd152: sin_out <= 13'b0100110001000;
                8'd153: sin_out <= 13'b0100101110100;
                8'd154: sin_out <= 13'b0100101011111;
                8'd155: sin_out <= 13'b0100101001011;
                8'd156: sin_out <= 13'b0100100110111;
                8'd157: sin_out <= 13'b0100100100010;
                8'd158: sin_out <= 13'b0100100001101;
                8'd159: sin_out <= 13'b0100011111000;
                8'd160: sin_out <= 13'b0100011100100;
                8'd161: sin_out <= 13'b0100011001111;
                8'd162: sin_out <= 13'b0100010111010;
                8'd163: sin_out <= 13'b0100010100101;
                8'd164: sin_out <= 13'b0100010001111;
                8'd165: sin_out <= 13'b0100001111010;
                8'd166: sin_out <= 13'b0100001100101;
                8'd167: sin_out <= 13'b0100001001111;
                8'd168: sin_out <= 13'b0100000111010;
                8'd169: sin_out <= 13'b0100000100100;
                8'd170: sin_out <= 13'b0100000001110;
                8'd171: sin_out <= 13'b0011111111001;
                8'd172: sin_out <= 13'b0011111100011;
                8'd173: sin_out <= 13'b0011111001101;
                8'd174: sin_out <= 13'b0011110110111;
                8'd175: sin_out <= 13'b0011110100001;
                8'd176: sin_out <= 13'b0011110001011;
                8'd177: sin_out <= 13'b0011101110101;
                8'd178: sin_out <= 13'b0011101011110;
                8'd179: sin_out <= 13'b0011101001000;
                8'd180: sin_out <= 13'b0011100110010;
                8'd181: sin_out <= 13'b0011100011011;
                8'd182: sin_out <= 13'b0011100000101;
                8'd183: sin_out <= 13'b0011011101110;
                8'd184: sin_out <= 13'b0011011010111;
                8'd185: sin_out <= 13'b0011011000001;
                8'd186: sin_out <= 13'b0011010101010;
                8'd187: sin_out <= 13'b0011010010011;
                8'd188: sin_out <= 13'b0011001111100;
                8'd189: sin_out <= 13'b0011001100101;
                8'd190: sin_out <= 13'b0011001001110;
                8'd191: sin_out <= 13'b0011000110111;
                8'd192: sin_out <= 13'b0011000011111;
                8'd193: sin_out <= 13'b0011000001000;
                8'd194: sin_out <= 13'b0010111110001;
                8'd195: sin_out <= 13'b0010111011010;
                8'd196: sin_out <= 13'b0010111000010;
                8'd197: sin_out <= 13'b0010110101011;
                8'd198: sin_out <= 13'b0010110010011;
                8'd199: sin_out <= 13'b0010101111100;
                8'd200: sin_out <= 13'b0010101100100;
                8'd201: sin_out <= 13'b0010101001100;
                8'd202: sin_out <= 13'b0010100110100;
                8'd203: sin_out <= 13'b0010100011101;
                8'd204: sin_out <= 13'b0010100000101;
                8'd205: sin_out <= 13'b0010011101101;
                8'd206: sin_out <= 13'b0010011010101;
                8'd207: sin_out <= 13'b0010010111101;
                8'd208: sin_out <= 13'b0010010100101;
                8'd209: sin_out <= 13'b0010010001101;
                8'd210: sin_out <= 13'b0010001110101;
                8'd211: sin_out <= 13'b0010001011101;
                8'd212: sin_out <= 13'b0010001000100;
                8'd213: sin_out <= 13'b0010000101100;
                8'd214: sin_out <= 13'b0010000010100;
                8'd215: sin_out <= 13'b0001111111100;
                8'd216: sin_out <= 13'b0001111100011;
                8'd217: sin_out <= 13'b0001111001011;
                8'd218: sin_out <= 13'b0001110110010;
                8'd219: sin_out <= 13'b0001110011010;
                8'd220: sin_out <= 13'b0001110000001;
                8'd221: sin_out <= 13'b0001101101001;
                8'd222: sin_out <= 13'b0001101010000;
                8'd223: sin_out <= 13'b0001100111000;
                8'd224: sin_out <= 13'b0001100011111;
                8'd225: sin_out <= 13'b0001100000110;
                8'd226: sin_out <= 13'b0001011101110;
                8'd227: sin_out <= 13'b0001011010101;
                8'd228: sin_out <= 13'b0001010111100;
                8'd229: sin_out <= 13'b0001010100011;
                8'd230: sin_out <= 13'b0001010001011;
                8'd231: sin_out <= 13'b0001001110010;
                8'd232: sin_out <= 13'b0001001011001;
                8'd233: sin_out <= 13'b0001001000000;
                8'd234: sin_out <= 13'b0001000100111;
                8'd235: sin_out <= 13'b0001000001110;
                8'd236: sin_out <= 13'b0000111110101;
                8'd237: sin_out <= 13'b0000111011100;
                8'd238: sin_out <= 13'b0000111000011;
                8'd239: sin_out <= 13'b0000110101010;
                8'd240: sin_out <= 13'b0000110010001;
                8'd241: sin_out <= 13'b0000101111000;
                8'd242: sin_out <= 13'b0000101011111;
                8'd243: sin_out <= 13'b0000101000110;
                8'd244: sin_out <= 13'b0000100101101;
                8'd245: sin_out <= 13'b0000100010100;
                8'd246: sin_out <= 13'b0000011111011;
                8'd247: sin_out <= 13'b0000011100010;
                8'd248: sin_out <= 13'b0000011001001;
                8'd249: sin_out <= 13'b0000010110000;
                8'd250: sin_out <= 13'b0000010010111;
                8'd251: sin_out <= 13'b0000001111110;
                8'd252: sin_out <= 13'b0000001100101;
                8'd253: sin_out <= 13'b0000001001011;
                8'd254: sin_out <= 13'b0000000110010;
                8'd255: sin_out <= 13'b0000000011001;
            endcase
        end
    endcase
end

endmodule
