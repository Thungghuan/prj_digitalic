module module_sin(sin_in, sin_out);

input [9:0] sin_in;
output [13:0] sin_out;

reg [13:0] out;

wire [1:0] high;
wire [7:0] low;

assign { high, low } = sin_in;

assign sin_out = out;

always @(*)
begin
    case (high)
        2'b00: 
        begin
            case (low)
                8'd000: out <= 14'b00000000000000;
                8'd001: out <= 14'b00000000011001;
                8'd002: out <= 14'b00000000110010;
                8'd003: out <= 14'b00000001001011;
                8'd004: out <= 14'b00000001100101;
                8'd005: out <= 14'b00000001111110;
                8'd006: out <= 14'b00000010010111;
                8'd007: out <= 14'b00000010110000;
                8'd008: out <= 14'b00000011001001;
                8'd009: out <= 14'b00000011100010;
                8'd010: out <= 14'b00000011111011;
                8'd011: out <= 14'b00000100010100;
                8'd012: out <= 14'b00000100101101;
                8'd013: out <= 14'b00000101000110;
                8'd014: out <= 14'b00000101011111;
                8'd015: out <= 14'b00000101111000;
                8'd016: out <= 14'b00000110010001;
                8'd017: out <= 14'b00000110101010;
                8'd018: out <= 14'b00000111000011;
                8'd019: out <= 14'b00000111011100;
                8'd020: out <= 14'b00000111110101;
                8'd021: out <= 14'b00001000001110;
                8'd022: out <= 14'b00001000100111;
                8'd023: out <= 14'b00001001000000;
                8'd024: out <= 14'b00001001011001;
                8'd025: out <= 14'b00001001110010;
                8'd026: out <= 14'b00001010001011;
                8'd027: out <= 14'b00001010100011;
                8'd028: out <= 14'b00001010111100;
                8'd029: out <= 14'b00001011010101;
                8'd030: out <= 14'b00001011101110;
                8'd031: out <= 14'b00001100000110;
                8'd032: out <= 14'b00001100011111;
                8'd033: out <= 14'b00001100111000;
                8'd034: out <= 14'b00001101010000;
                8'd035: out <= 14'b00001101101001;
                8'd036: out <= 14'b00001110000001;
                8'd037: out <= 14'b00001110011010;
                8'd038: out <= 14'b00001110110010;
                8'd039: out <= 14'b00001111001011;
                8'd040: out <= 14'b00001111100011;
                8'd041: out <= 14'b00001111111100;
                8'd042: out <= 14'b00010000010100;
                8'd043: out <= 14'b00010000101100;
                8'd044: out <= 14'b00010001000100;
                8'd045: out <= 14'b00010001011101;
                8'd046: out <= 14'b00010001110101;
                8'd047: out <= 14'b00010010001101;
                8'd048: out <= 14'b00010010100101;
                8'd049: out <= 14'b00010010111101;
                8'd050: out <= 14'b00010011010101;
                8'd051: out <= 14'b00010011101101;
                8'd052: out <= 14'b00010100000101;
                8'd053: out <= 14'b00010100011101;
                8'd054: out <= 14'b00010100110100;
                8'd055: out <= 14'b00010101001100;
                8'd056: out <= 14'b00010101100100;
                8'd057: out <= 14'b00010101111100;
                8'd058: out <= 14'b00010110010011;
                8'd059: out <= 14'b00010110101011;
                8'd060: out <= 14'b00010111000010;
                8'd061: out <= 14'b00010111011010;
                8'd062: out <= 14'b00010111110001;
                8'd063: out <= 14'b00011000001000;
                8'd064: out <= 14'b00011000011111;
                8'd065: out <= 14'b00011000110111;
                8'd066: out <= 14'b00011001001110;
                8'd067: out <= 14'b00011001100101;
                8'd068: out <= 14'b00011001111100;
                8'd069: out <= 14'b00011010010011;
                8'd070: out <= 14'b00011010101010;
                8'd071: out <= 14'b00011011000001;
                8'd072: out <= 14'b00011011010111;
                8'd073: out <= 14'b00011011101110;
                8'd074: out <= 14'b00011100000101;
                8'd075: out <= 14'b00011100011011;
                8'd076: out <= 14'b00011100110010;
                8'd077: out <= 14'b00011101001000;
                8'd078: out <= 14'b00011101011110;
                8'd079: out <= 14'b00011101110101;
                8'd080: out <= 14'b00011110001011;
                8'd081: out <= 14'b00011110100001;
                8'd082: out <= 14'b00011110110111;
                8'd083: out <= 14'b00011111001101;
                8'd084: out <= 14'b00011111100011;
                8'd085: out <= 14'b00011111111001;
                8'd086: out <= 14'b00100000001110;
                8'd087: out <= 14'b00100000100100;
                8'd088: out <= 14'b00100000111010;
                8'd089: out <= 14'b00100001001111;
                8'd090: out <= 14'b00100001100101;
                8'd091: out <= 14'b00100001111010;
                8'd092: out <= 14'b00100010001111;
                8'd093: out <= 14'b00100010100101;
                8'd094: out <= 14'b00100010111010;
                8'd095: out <= 14'b00100011001111;
                8'd096: out <= 14'b00100011100100;
                8'd097: out <= 14'b00100011111000;
                8'd098: out <= 14'b00100100001101;
                8'd099: out <= 14'b00100100100010;
                8'd100: out <= 14'b00100100110111;
                8'd101: out <= 14'b00100101001011;
                8'd102: out <= 14'b00100101011111;
                8'd103: out <= 14'b00100101110100;
                8'd104: out <= 14'b00100110001000;
                8'd105: out <= 14'b00100110011100;
                8'd106: out <= 14'b00100110110000;
                8'd107: out <= 14'b00100111000100;
                8'd108: out <= 14'b00100111011000;
                8'd109: out <= 14'b00100111101100;
                8'd110: out <= 14'b00100111111111;
                8'd111: out <= 14'b00101000010011;
                8'd112: out <= 14'b00101000100110;
                8'd113: out <= 14'b00101000111010;
                8'd114: out <= 14'b00101001001101;
                8'd115: out <= 14'b00101001100000;
                8'd116: out <= 14'b00101001110011;
                8'd117: out <= 14'b00101010000110;
                8'd118: out <= 14'b00101010011001;
                8'd119: out <= 14'b00101010101100;
                8'd120: out <= 14'b00101010111111;
                8'd121: out <= 14'b00101011010001;
                8'd122: out <= 14'b00101011100100;
                8'd123: out <= 14'b00101011110110;
                8'd124: out <= 14'b00101100001000;
                8'd125: out <= 14'b00101100011011;
                8'd126: out <= 14'b00101100101101;
                8'd127: out <= 14'b00101100111110;
                8'd128: out <= 14'b00101101010000;
                8'd129: out <= 14'b00101101100010;
                8'd130: out <= 14'b00101101110100;
                8'd131: out <= 14'b00101110000101;
                8'd132: out <= 14'b00101110010111;
                8'd133: out <= 14'b00101110101000;
                8'd134: out <= 14'b00101110111001;
                8'd135: out <= 14'b00101111001010;
                8'd136: out <= 14'b00101111011011;
                8'd137: out <= 14'b00101111101100;
                8'd138: out <= 14'b00101111111100;
                8'd139: out <= 14'b00110000001101;
                8'd140: out <= 14'b00110000011110;
                8'd141: out <= 14'b00110000101110;
                8'd142: out <= 14'b00110000111110;
                8'd143: out <= 14'b00110001001110;
                8'd144: out <= 14'b00110001011110;
                8'd145: out <= 14'b00110001101110;
                8'd146: out <= 14'b00110001111110;
                8'd147: out <= 14'b00110010001110;
                8'd148: out <= 14'b00110010011101;
                8'd149: out <= 14'b00110010101100;
                8'd150: out <= 14'b00110010111100;
                8'd151: out <= 14'b00110011001011;
                8'd152: out <= 14'b00110011011010;
                8'd153: out <= 14'b00110011101001;
                8'd154: out <= 14'b00110011111000;
                8'd155: out <= 14'b00110100000110;
                8'd156: out <= 14'b00110100010101;
                8'd157: out <= 14'b00110100100011;
                8'd158: out <= 14'b00110100110010;
                8'd159: out <= 14'b00110101000000;
                8'd160: out <= 14'b00110101001110;
                8'd161: out <= 14'b00110101011100;
                8'd162: out <= 14'b00110101101001;
                8'd163: out <= 14'b00110101110111;
                8'd164: out <= 14'b00110110000101;
                8'd165: out <= 14'b00110110010010;
                8'd166: out <= 14'b00110110011111;
                8'd167: out <= 14'b00110110101100;
                8'd168: out <= 14'b00110110111001;
                8'd169: out <= 14'b00110111000110;
                8'd170: out <= 14'b00110111010011;
                8'd171: out <= 14'b00110111011111;
                8'd172: out <= 14'b00110111101100;
                8'd173: out <= 14'b00110111111000;
                8'd174: out <= 14'b00111000000100;
                8'd175: out <= 14'b00111000010000;
                8'd176: out <= 14'b00111000011100;
                8'd177: out <= 14'b00111000101000;
                8'd178: out <= 14'b00111000110100;
                8'd179: out <= 14'b00111000111111;
                8'd180: out <= 14'b00111001001011;
                8'd181: out <= 14'b00111001010110;
                8'd182: out <= 14'b00111001100001;
                8'd183: out <= 14'b00111001101100;
                8'd184: out <= 14'b00111001110111;
                8'd185: out <= 14'b00111010000001;
                8'd186: out <= 14'b00111010001100;
                8'd187: out <= 14'b00111010010110;
                8'd188: out <= 14'b00111010100001;
                8'd189: out <= 14'b00111010101011;
                8'd190: out <= 14'b00111010110101;
                8'd191: out <= 14'b00111010111111;
                8'd192: out <= 14'b00111011001000;
                8'd193: out <= 14'b00111011010010;
                8'd194: out <= 14'b00111011011011;
                8'd195: out <= 14'b00111011100100;
                8'd196: out <= 14'b00111011101110;
                8'd197: out <= 14'b00111011110111;
                8'd198: out <= 14'b00111011111111;
                8'd199: out <= 14'b00111100001000;
                8'd200: out <= 14'b00111100010001;
                8'd201: out <= 14'b00111100011001;
                8'd202: out <= 14'b00111100100001;
                8'd203: out <= 14'b00111100101001;
                8'd204: out <= 14'b00111100110001;
                8'd205: out <= 14'b00111100111001;
                8'd206: out <= 14'b00111101000001;
                8'd207: out <= 14'b00111101001000;
                8'd208: out <= 14'b00111101010000;
                8'd209: out <= 14'b00111101010111;
                8'd210: out <= 14'b00111101011110;
                8'd211: out <= 14'b00111101100101;
                8'd212: out <= 14'b00111101101100;
                8'd213: out <= 14'b00111101110010;
                8'd214: out <= 14'b00111101111001;
                8'd215: out <= 14'b00111101111111;
                8'd216: out <= 14'b00111110000101;
                8'd217: out <= 14'b00111110001011;
                8'd218: out <= 14'b00111110010001;
                8'd219: out <= 14'b00111110010111;
                8'd220: out <= 14'b00111110011100;
                8'd221: out <= 14'b00111110100010;
                8'd222: out <= 14'b00111110100111;
                8'd223: out <= 14'b00111110101100;
                8'd224: out <= 14'b00111110110001;
                8'd225: out <= 14'b00111110110110;
                8'd226: out <= 14'b00111110111011;
                8'd227: out <= 14'b00111110111111;
                8'd228: out <= 14'b00111111000100;
                8'd229: out <= 14'b00111111001000;
                8'd230: out <= 14'b00111111001100;
                8'd231: out <= 14'b00111111010000;
                8'd232: out <= 14'b00111111010100;
                8'd233: out <= 14'b00111111010111;
                8'd234: out <= 14'b00111111011011;
                8'd235: out <= 14'b00111111011110;
                8'd236: out <= 14'b00111111100001;
                8'd237: out <= 14'b00111111100100;
                8'd238: out <= 14'b00111111100111;
                8'd239: out <= 14'b00111111101010;
                8'd240: out <= 14'b00111111101100;
                8'd241: out <= 14'b00111111101111;
                8'd242: out <= 14'b00111111110001;
                8'd243: out <= 14'b00111111110011;
                8'd244: out <= 14'b00111111110101;
                8'd245: out <= 14'b00111111110111;
                8'd246: out <= 14'b00111111111000;
                8'd247: out <= 14'b00111111111010;
                8'd248: out <= 14'b00111111111011;
                8'd249: out <= 14'b00111111111100;
                8'd250: out <= 14'b00111111111101;
                8'd251: out <= 14'b00111111111110;
                8'd252: out <= 14'b00111111111111;
                8'd253: out <= 14'b00111111111111;
                8'd254: out <= 14'b01000000000000;
                8'd255: out <= 14'b01000000000000;
            endcase        end
        2'b01: 
        begin
            case (low)
                8'd000: out <= 14'b01000000000000;
                8'd001: out <= 14'b01000000000000;
                8'd002: out <= 14'b01000000000000;
                8'd003: out <= 14'b00111111111111;
                8'd004: out <= 14'b00111111111111;
                8'd005: out <= 14'b00111111111110;
                8'd006: out <= 14'b00111111111101;
                8'd007: out <= 14'b00111111111100;
                8'd008: out <= 14'b00111111111011;
                8'd009: out <= 14'b00111111111010;
                8'd010: out <= 14'b00111111111000;
                8'd011: out <= 14'b00111111110111;
                8'd012: out <= 14'b00111111110101;
                8'd013: out <= 14'b00111111110011;
                8'd014: out <= 14'b00111111110001;
                8'd015: out <= 14'b00111111101111;
                8'd016: out <= 14'b00111111101100;
                8'd017: out <= 14'b00111111101010;
                8'd018: out <= 14'b00111111100111;
                8'd019: out <= 14'b00111111100100;
                8'd020: out <= 14'b00111111100001;
                8'd021: out <= 14'b00111111011110;
                8'd022: out <= 14'b00111111011011;
                8'd023: out <= 14'b00111111010111;
                8'd024: out <= 14'b00111111010100;
                8'd025: out <= 14'b00111111010000;
                8'd026: out <= 14'b00111111001100;
                8'd027: out <= 14'b00111111001000;
                8'd028: out <= 14'b00111111000100;
                8'd029: out <= 14'b00111110111111;
                8'd030: out <= 14'b00111110111011;
                8'd031: out <= 14'b00111110110110;
                8'd032: out <= 14'b00111110110001;
                8'd033: out <= 14'b00111110101100;
                8'd034: out <= 14'b00111110100111;
                8'd035: out <= 14'b00111110100010;
                8'd036: out <= 14'b00111110011100;
                8'd037: out <= 14'b00111110010111;
                8'd038: out <= 14'b00111110010001;
                8'd039: out <= 14'b00111110001011;
                8'd040: out <= 14'b00111110000101;
                8'd041: out <= 14'b00111101111111;
                8'd042: out <= 14'b00111101111001;
                8'd043: out <= 14'b00111101110010;
                8'd044: out <= 14'b00111101101100;
                8'd045: out <= 14'b00111101100101;
                8'd046: out <= 14'b00111101011110;
                8'd047: out <= 14'b00111101010111;
                8'd048: out <= 14'b00111101010000;
                8'd049: out <= 14'b00111101001000;
                8'd050: out <= 14'b00111101000001;
                8'd051: out <= 14'b00111100111001;
                8'd052: out <= 14'b00111100110001;
                8'd053: out <= 14'b00111100101001;
                8'd054: out <= 14'b00111100100001;
                8'd055: out <= 14'b00111100011001;
                8'd056: out <= 14'b00111100010001;
                8'd057: out <= 14'b00111100001000;
                8'd058: out <= 14'b00111011111111;
                8'd059: out <= 14'b00111011110111;
                8'd060: out <= 14'b00111011101110;
                8'd061: out <= 14'b00111011100100;
                8'd062: out <= 14'b00111011011011;
                8'd063: out <= 14'b00111011010010;
                8'd064: out <= 14'b00111011001000;
                8'd065: out <= 14'b00111010111111;
                8'd066: out <= 14'b00111010110101;
                8'd067: out <= 14'b00111010101011;
                8'd068: out <= 14'b00111010100001;
                8'd069: out <= 14'b00111010010110;
                8'd070: out <= 14'b00111010001100;
                8'd071: out <= 14'b00111010000001;
                8'd072: out <= 14'b00111001110111;
                8'd073: out <= 14'b00111001101100;
                8'd074: out <= 14'b00111001100001;
                8'd075: out <= 14'b00111001010110;
                8'd076: out <= 14'b00111001001011;
                8'd077: out <= 14'b00111000111111;
                8'd078: out <= 14'b00111000110100;
                8'd079: out <= 14'b00111000101000;
                8'd080: out <= 14'b00111000011100;
                8'd081: out <= 14'b00111000010000;
                8'd082: out <= 14'b00111000000100;
                8'd083: out <= 14'b00110111111000;
                8'd084: out <= 14'b00110111101100;
                8'd085: out <= 14'b00110111011111;
                8'd086: out <= 14'b00110111010011;
                8'd087: out <= 14'b00110111000110;
                8'd088: out <= 14'b00110110111001;
                8'd089: out <= 14'b00110110101100;
                8'd090: out <= 14'b00110110011111;
                8'd091: out <= 14'b00110110010010;
                8'd092: out <= 14'b00110110000101;
                8'd093: out <= 14'b00110101110111;
                8'd094: out <= 14'b00110101101001;
                8'd095: out <= 14'b00110101011100;
                8'd096: out <= 14'b00110101001110;
                8'd097: out <= 14'b00110101000000;
                8'd098: out <= 14'b00110100110010;
                8'd099: out <= 14'b00110100100011;
                8'd100: out <= 14'b00110100010101;
                8'd101: out <= 14'b00110100000110;
                8'd102: out <= 14'b00110011111000;
                8'd103: out <= 14'b00110011101001;
                8'd104: out <= 14'b00110011011010;
                8'd105: out <= 14'b00110011001011;
                8'd106: out <= 14'b00110010111100;
                8'd107: out <= 14'b00110010101100;
                8'd108: out <= 14'b00110010011101;
                8'd109: out <= 14'b00110010001110;
                8'd110: out <= 14'b00110001111110;
                8'd111: out <= 14'b00110001101110;
                8'd112: out <= 14'b00110001011110;
                8'd113: out <= 14'b00110001001110;
                8'd114: out <= 14'b00110000111110;
                8'd115: out <= 14'b00110000101110;
                8'd116: out <= 14'b00110000011110;
                8'd117: out <= 14'b00110000001101;
                8'd118: out <= 14'b00101111111100;
                8'd119: out <= 14'b00101111101100;
                8'd120: out <= 14'b00101111011011;
                8'd121: out <= 14'b00101111001010;
                8'd122: out <= 14'b00101110111001;
                8'd123: out <= 14'b00101110101000;
                8'd124: out <= 14'b00101110010111;
                8'd125: out <= 14'b00101110000101;
                8'd126: out <= 14'b00101101110100;
                8'd127: out <= 14'b00101101100010;
                8'd128: out <= 14'b00101101010000;
                8'd129: out <= 14'b00101100111110;
                8'd130: out <= 14'b00101100101101;
                8'd131: out <= 14'b00101100011011;
                8'd132: out <= 14'b00101100001000;
                8'd133: out <= 14'b00101011110110;
                8'd134: out <= 14'b00101011100100;
                8'd135: out <= 14'b00101011010001;
                8'd136: out <= 14'b00101010111111;
                8'd137: out <= 14'b00101010101100;
                8'd138: out <= 14'b00101010011001;
                8'd139: out <= 14'b00101010000110;
                8'd140: out <= 14'b00101001110011;
                8'd141: out <= 14'b00101001100000;
                8'd142: out <= 14'b00101001001101;
                8'd143: out <= 14'b00101000111010;
                8'd144: out <= 14'b00101000100110;
                8'd145: out <= 14'b00101000010011;
                8'd146: out <= 14'b00100111111111;
                8'd147: out <= 14'b00100111101100;
                8'd148: out <= 14'b00100111011000;
                8'd149: out <= 14'b00100111000100;
                8'd150: out <= 14'b00100110110000;
                8'd151: out <= 14'b00100110011100;
                8'd152: out <= 14'b00100110001000;
                8'd153: out <= 14'b00100101110100;
                8'd154: out <= 14'b00100101011111;
                8'd155: out <= 14'b00100101001011;
                8'd156: out <= 14'b00100100110111;
                8'd157: out <= 14'b00100100100010;
                8'd158: out <= 14'b00100100001101;
                8'd159: out <= 14'b00100011111000;
                8'd160: out <= 14'b00100011100100;
                8'd161: out <= 14'b00100011001111;
                8'd162: out <= 14'b00100010111010;
                8'd163: out <= 14'b00100010100101;
                8'd164: out <= 14'b00100010001111;
                8'd165: out <= 14'b00100001111010;
                8'd166: out <= 14'b00100001100101;
                8'd167: out <= 14'b00100001001111;
                8'd168: out <= 14'b00100000111010;
                8'd169: out <= 14'b00100000100100;
                8'd170: out <= 14'b00100000001110;
                8'd171: out <= 14'b00011111111001;
                8'd172: out <= 14'b00011111100011;
                8'd173: out <= 14'b00011111001101;
                8'd174: out <= 14'b00011110110111;
                8'd175: out <= 14'b00011110100001;
                8'd176: out <= 14'b00011110001011;
                8'd177: out <= 14'b00011101110101;
                8'd178: out <= 14'b00011101011110;
                8'd179: out <= 14'b00011101001000;
                8'd180: out <= 14'b00011100110010;
                8'd181: out <= 14'b00011100011011;
                8'd182: out <= 14'b00011100000101;
                8'd183: out <= 14'b00011011101110;
                8'd184: out <= 14'b00011011010111;
                8'd185: out <= 14'b00011011000001;
                8'd186: out <= 14'b00011010101010;
                8'd187: out <= 14'b00011010010011;
                8'd188: out <= 14'b00011001111100;
                8'd189: out <= 14'b00011001100101;
                8'd190: out <= 14'b00011001001110;
                8'd191: out <= 14'b00011000110111;
                8'd192: out <= 14'b00011000011111;
                8'd193: out <= 14'b00011000001000;
                8'd194: out <= 14'b00010111110001;
                8'd195: out <= 14'b00010111011010;
                8'd196: out <= 14'b00010111000010;
                8'd197: out <= 14'b00010110101011;
                8'd198: out <= 14'b00010110010011;
                8'd199: out <= 14'b00010101111100;
                8'd200: out <= 14'b00010101100100;
                8'd201: out <= 14'b00010101001100;
                8'd202: out <= 14'b00010100110100;
                8'd203: out <= 14'b00010100011101;
                8'd204: out <= 14'b00010100000101;
                8'd205: out <= 14'b00010011101101;
                8'd206: out <= 14'b00010011010101;
                8'd207: out <= 14'b00010010111101;
                8'd208: out <= 14'b00010010100101;
                8'd209: out <= 14'b00010010001101;
                8'd210: out <= 14'b00010001110101;
                8'd211: out <= 14'b00010001011101;
                8'd212: out <= 14'b00010001000100;
                8'd213: out <= 14'b00010000101100;
                8'd214: out <= 14'b00010000010100;
                8'd215: out <= 14'b00001111111100;
                8'd216: out <= 14'b00001111100011;
                8'd217: out <= 14'b00001111001011;
                8'd218: out <= 14'b00001110110010;
                8'd219: out <= 14'b00001110011010;
                8'd220: out <= 14'b00001110000001;
                8'd221: out <= 14'b00001101101001;
                8'd222: out <= 14'b00001101010000;
                8'd223: out <= 14'b00001100111000;
                8'd224: out <= 14'b00001100011111;
                8'd225: out <= 14'b00001100000110;
                8'd226: out <= 14'b00001011101110;
                8'd227: out <= 14'b00001011010101;
                8'd228: out <= 14'b00001010111100;
                8'd229: out <= 14'b00001010100011;
                8'd230: out <= 14'b00001010001011;
                8'd231: out <= 14'b00001001110010;
                8'd232: out <= 14'b00001001011001;
                8'd233: out <= 14'b00001001000000;
                8'd234: out <= 14'b00001000100111;
                8'd235: out <= 14'b00001000001110;
                8'd236: out <= 14'b00000111110101;
                8'd237: out <= 14'b00000111011100;
                8'd238: out <= 14'b00000111000011;
                8'd239: out <= 14'b00000110101010;
                8'd240: out <= 14'b00000110010001;
                8'd241: out <= 14'b00000101111000;
                8'd242: out <= 14'b00000101011111;
                8'd243: out <= 14'b00000101000110;
                8'd244: out <= 14'b00000100101101;
                8'd245: out <= 14'b00000100010100;
                8'd246: out <= 14'b00000011111011;
                8'd247: out <= 14'b00000011100010;
                8'd248: out <= 14'b00000011001001;
                8'd249: out <= 14'b00000010110000;
                8'd250: out <= 14'b00000010010111;
                8'd251: out <= 14'b00000001111110;
                8'd252: out <= 14'b00000001100101;
                8'd253: out <= 14'b00000001001011;
                8'd254: out <= 14'b00000000110010;
                8'd255: out <= 14'b00000000011001;
            endcase        end
        2'b10: 
        begin
            case (low)
                8'd000: out <= 14'b00000000000000;
                8'd001: out <= 14'b11111111100111;
                8'd002: out <= 14'b11111111001110;
                8'd003: out <= 14'b11111110110101;
                8'd004: out <= 14'b11111110011011;
                8'd005: out <= 14'b11111110000010;
                8'd006: out <= 14'b11111101101001;
                8'd007: out <= 14'b11111101010000;
                8'd008: out <= 14'b11111100110111;
                8'd009: out <= 14'b11111100011110;
                8'd010: out <= 14'b11111100000101;
                8'd011: out <= 14'b11111011101100;
                8'd012: out <= 14'b11111011010011;
                8'd013: out <= 14'b11111010111010;
                8'd014: out <= 14'b11111010100001;
                8'd015: out <= 14'b11111010001000;
                8'd016: out <= 14'b11111001101111;
                8'd017: out <= 14'b11111001010110;
                8'd018: out <= 14'b11111000111101;
                8'd019: out <= 14'b11111000100100;
                8'd020: out <= 14'b11111000001011;
                8'd021: out <= 14'b11110111110010;
                8'd022: out <= 14'b11110111011001;
                8'd023: out <= 14'b11110111000000;
                8'd024: out <= 14'b11110110100111;
                8'd025: out <= 14'b11110110001110;
                8'd026: out <= 14'b11110101110101;
                8'd027: out <= 14'b11110101011101;
                8'd028: out <= 14'b11110101000100;
                8'd029: out <= 14'b11110100101011;
                8'd030: out <= 14'b11110100010010;
                8'd031: out <= 14'b11110011111010;
                8'd032: out <= 14'b11110011100001;
                8'd033: out <= 14'b11110011001000;
                8'd034: out <= 14'b11110010110000;
                8'd035: out <= 14'b11110010010111;
                8'd036: out <= 14'b11110001111111;
                8'd037: out <= 14'b11110001100110;
                8'd038: out <= 14'b11110001001110;
                8'd039: out <= 14'b11110000110101;
                8'd040: out <= 14'b11110000011101;
                8'd041: out <= 14'b11110000000100;
                8'd042: out <= 14'b11101111101100;
                8'd043: out <= 14'b11101111010100;
                8'd044: out <= 14'b11101110111100;
                8'd045: out <= 14'b11101110100011;
                8'd046: out <= 14'b11101110001011;
                8'd047: out <= 14'b11101101110011;
                8'd048: out <= 14'b11101101011011;
                8'd049: out <= 14'b11101101000011;
                8'd050: out <= 14'b11101100101011;
                8'd051: out <= 14'b11101100010011;
                8'd052: out <= 14'b11101011111011;
                8'd053: out <= 14'b11101011100011;
                8'd054: out <= 14'b11101011001100;
                8'd055: out <= 14'b11101010110100;
                8'd056: out <= 14'b11101010011100;
                8'd057: out <= 14'b11101010000100;
                8'd058: out <= 14'b11101001101101;
                8'd059: out <= 14'b11101001010101;
                8'd060: out <= 14'b11101000111110;
                8'd061: out <= 14'b11101000100110;
                8'd062: out <= 14'b11101000001111;
                8'd063: out <= 14'b11100111111000;
                8'd064: out <= 14'b11100111100001;
                8'd065: out <= 14'b11100111001001;
                8'd066: out <= 14'b11100110110010;
                8'd067: out <= 14'b11100110011011;
                8'd068: out <= 14'b11100110000100;
                8'd069: out <= 14'b11100101101101;
                8'd070: out <= 14'b11100101010110;
                8'd071: out <= 14'b11100100111111;
                8'd072: out <= 14'b11100100101001;
                8'd073: out <= 14'b11100100010010;
                8'd074: out <= 14'b11100011111011;
                8'd075: out <= 14'b11100011100101;
                8'd076: out <= 14'b11100011001110;
                8'd077: out <= 14'b11100010111000;
                8'd078: out <= 14'b11100010100010;
                8'd079: out <= 14'b11100010001011;
                8'd080: out <= 14'b11100001110101;
                8'd081: out <= 14'b11100001011111;
                8'd082: out <= 14'b11100001001001;
                8'd083: out <= 14'b11100000110011;
                8'd084: out <= 14'b11100000011101;
                8'd085: out <= 14'b11100000000111;
                8'd086: out <= 14'b11011111110010;
                8'd087: out <= 14'b11011111011100;
                8'd088: out <= 14'b11011111000110;
                8'd089: out <= 14'b11011110110001;
                8'd090: out <= 14'b11011110011011;
                8'd091: out <= 14'b11011110000110;
                8'd092: out <= 14'b11011101110001;
                8'd093: out <= 14'b11011101011011;
                8'd094: out <= 14'b11011101000110;
                8'd095: out <= 14'b11011100110001;
                8'd096: out <= 14'b11011100011100;
                8'd097: out <= 14'b11011100001000;
                8'd098: out <= 14'b11011011110011;
                8'd099: out <= 14'b11011011011110;
                8'd100: out <= 14'b11011011001001;
                8'd101: out <= 14'b11011010110101;
                8'd102: out <= 14'b11011010100001;
                8'd103: out <= 14'b11011010001100;
                8'd104: out <= 14'b11011001111000;
                8'd105: out <= 14'b11011001100100;
                8'd106: out <= 14'b11011001010000;
                8'd107: out <= 14'b11011000111100;
                8'd108: out <= 14'b11011000101000;
                8'd109: out <= 14'b11011000010100;
                8'd110: out <= 14'b11011000000001;
                8'd111: out <= 14'b11010111101101;
                8'd112: out <= 14'b11010111011010;
                8'd113: out <= 14'b11010111000110;
                8'd114: out <= 14'b11010110110011;
                8'd115: out <= 14'b11010110100000;
                8'd116: out <= 14'b11010110001101;
                8'd117: out <= 14'b11010101111010;
                8'd118: out <= 14'b11010101100111;
                8'd119: out <= 14'b11010101010100;
                8'd120: out <= 14'b11010101000001;
                8'd121: out <= 14'b11010100101111;
                8'd122: out <= 14'b11010100011100;
                8'd123: out <= 14'b11010100001010;
                8'd124: out <= 14'b11010011111000;
                8'd125: out <= 14'b11010011100101;
                8'd126: out <= 14'b11010011010011;
                8'd127: out <= 14'b11010011000010;
                8'd128: out <= 14'b11010010110000;
                8'd129: out <= 14'b11010010011110;
                8'd130: out <= 14'b11010010001100;
                8'd131: out <= 14'b11010001111011;
                8'd132: out <= 14'b11010001101001;
                8'd133: out <= 14'b11010001011000;
                8'd134: out <= 14'b11010001000111;
                8'd135: out <= 14'b11010000110110;
                8'd136: out <= 14'b11010000100101;
                8'd137: out <= 14'b11010000010100;
                8'd138: out <= 14'b11010000000100;
                8'd139: out <= 14'b11001111110011;
                8'd140: out <= 14'b11001111100010;
                8'd141: out <= 14'b11001111010010;
                8'd142: out <= 14'b11001111000010;
                8'd143: out <= 14'b11001110110010;
                8'd144: out <= 14'b11001110100010;
                8'd145: out <= 14'b11001110010010;
                8'd146: out <= 14'b11001110000010;
                8'd147: out <= 14'b11001101110010;
                8'd148: out <= 14'b11001101100011;
                8'd149: out <= 14'b11001101010100;
                8'd150: out <= 14'b11001101000100;
                8'd151: out <= 14'b11001100110101;
                8'd152: out <= 14'b11001100100110;
                8'd153: out <= 14'b11001100010111;
                8'd154: out <= 14'b11001100001000;
                8'd155: out <= 14'b11001011111010;
                8'd156: out <= 14'b11001011101011;
                8'd157: out <= 14'b11001011011101;
                8'd158: out <= 14'b11001011001110;
                8'd159: out <= 14'b11001011000000;
                8'd160: out <= 14'b11001010110010;
                8'd161: out <= 14'b11001010100100;
                8'd162: out <= 14'b11001010010111;
                8'd163: out <= 14'b11001010001001;
                8'd164: out <= 14'b11001001111011;
                8'd165: out <= 14'b11001001101110;
                8'd166: out <= 14'b11001001100001;
                8'd167: out <= 14'b11001001010100;
                8'd168: out <= 14'b11001001000111;
                8'd169: out <= 14'b11001000111010;
                8'd170: out <= 14'b11001000101101;
                8'd171: out <= 14'b11001000100001;
                8'd172: out <= 14'b11001000010100;
                8'd173: out <= 14'b11001000001000;
                8'd174: out <= 14'b11000111111100;
                8'd175: out <= 14'b11000111110000;
                8'd176: out <= 14'b11000111100100;
                8'd177: out <= 14'b11000111011000;
                8'd178: out <= 14'b11000111001100;
                8'd179: out <= 14'b11000111000001;
                8'd180: out <= 14'b11000110110101;
                8'd181: out <= 14'b11000110101010;
                8'd182: out <= 14'b11000110011111;
                8'd183: out <= 14'b11000110010100;
                8'd184: out <= 14'b11000110001001;
                8'd185: out <= 14'b11000101111111;
                8'd186: out <= 14'b11000101110100;
                8'd187: out <= 14'b11000101101010;
                8'd188: out <= 14'b11000101011111;
                8'd189: out <= 14'b11000101010101;
                8'd190: out <= 14'b11000101001011;
                8'd191: out <= 14'b11000101000001;
                8'd192: out <= 14'b11000100111000;
                8'd193: out <= 14'b11000100101110;
                8'd194: out <= 14'b11000100100101;
                8'd195: out <= 14'b11000100011100;
                8'd196: out <= 14'b11000100010010;
                8'd197: out <= 14'b11000100001001;
                8'd198: out <= 14'b11000100000001;
                8'd199: out <= 14'b11000011111000;
                8'd200: out <= 14'b11000011101111;
                8'd201: out <= 14'b11000011100111;
                8'd202: out <= 14'b11000011011111;
                8'd203: out <= 14'b11000011010111;
                8'd204: out <= 14'b11000011001111;
                8'd205: out <= 14'b11000011000111;
                8'd206: out <= 14'b11000010111111;
                8'd207: out <= 14'b11000010111000;
                8'd208: out <= 14'b11000010110000;
                8'd209: out <= 14'b11000010101001;
                8'd210: out <= 14'b11000010100010;
                8'd211: out <= 14'b11000010011011;
                8'd212: out <= 14'b11000010010100;
                8'd213: out <= 14'b11000010001110;
                8'd214: out <= 14'b11000010000111;
                8'd215: out <= 14'b11000010000001;
                8'd216: out <= 14'b11000001111011;
                8'd217: out <= 14'b11000001110101;
                8'd218: out <= 14'b11000001101111;
                8'd219: out <= 14'b11000001101001;
                8'd220: out <= 14'b11000001100100;
                8'd221: out <= 14'b11000001011110;
                8'd222: out <= 14'b11000001011001;
                8'd223: out <= 14'b11000001010100;
                8'd224: out <= 14'b11000001001111;
                8'd225: out <= 14'b11000001001010;
                8'd226: out <= 14'b11000001000101;
                8'd227: out <= 14'b11000001000001;
                8'd228: out <= 14'b11000000111100;
                8'd229: out <= 14'b11000000111000;
                8'd230: out <= 14'b11000000110100;
                8'd231: out <= 14'b11000000110000;
                8'd232: out <= 14'b11000000101100;
                8'd233: out <= 14'b11000000101001;
                8'd234: out <= 14'b11000000100101;
                8'd235: out <= 14'b11000000100010;
                8'd236: out <= 14'b11000000011111;
                8'd237: out <= 14'b11000000011100;
                8'd238: out <= 14'b11000000011001;
                8'd239: out <= 14'b11000000010110;
                8'd240: out <= 14'b11000000010100;
                8'd241: out <= 14'b11000000010001;
                8'd242: out <= 14'b11000000001111;
                8'd243: out <= 14'b11000000001101;
                8'd244: out <= 14'b11000000001011;
                8'd245: out <= 14'b11000000001001;
                8'd246: out <= 14'b11000000001000;
                8'd247: out <= 14'b11000000000110;
                8'd248: out <= 14'b11000000000101;
                8'd249: out <= 14'b11000000000100;
                8'd250: out <= 14'b11000000000011;
                8'd251: out <= 14'b11000000000010;
                8'd252: out <= 14'b11000000000001;
                8'd253: out <= 14'b11000000000001;
                8'd254: out <= 14'b11000000000000;
                8'd255: out <= 14'b11000000000000;
            endcase        end
        2'b11: 
        begin
            case (low)
                8'd000: out <= 14'b11000000000000;
                8'd001: out <= 14'b11000000000000;
                8'd002: out <= 14'b11000000000000;
                8'd003: out <= 14'b11000000000001;
                8'd004: out <= 14'b11000000000001;
                8'd005: out <= 14'b11000000000010;
                8'd006: out <= 14'b11000000000011;
                8'd007: out <= 14'b11000000000100;
                8'd008: out <= 14'b11000000000101;
                8'd009: out <= 14'b11000000000110;
                8'd010: out <= 14'b11000000001000;
                8'd011: out <= 14'b11000000001001;
                8'd012: out <= 14'b11000000001011;
                8'd013: out <= 14'b11000000001101;
                8'd014: out <= 14'b11000000001111;
                8'd015: out <= 14'b11000000010001;
                8'd016: out <= 14'b11000000010100;
                8'd017: out <= 14'b11000000010110;
                8'd018: out <= 14'b11000000011001;
                8'd019: out <= 14'b11000000011100;
                8'd020: out <= 14'b11000000011111;
                8'd021: out <= 14'b11000000100010;
                8'd022: out <= 14'b11000000100101;
                8'd023: out <= 14'b11000000101001;
                8'd024: out <= 14'b11000000101100;
                8'd025: out <= 14'b11000000110000;
                8'd026: out <= 14'b11000000110100;
                8'd027: out <= 14'b11000000111000;
                8'd028: out <= 14'b11000000111100;
                8'd029: out <= 14'b11000001000001;
                8'd030: out <= 14'b11000001000101;
                8'd031: out <= 14'b11000001001010;
                8'd032: out <= 14'b11000001001111;
                8'd033: out <= 14'b11000001010100;
                8'd034: out <= 14'b11000001011001;
                8'd035: out <= 14'b11000001011110;
                8'd036: out <= 14'b11000001100100;
                8'd037: out <= 14'b11000001101001;
                8'd038: out <= 14'b11000001101111;
                8'd039: out <= 14'b11000001110101;
                8'd040: out <= 14'b11000001111011;
                8'd041: out <= 14'b11000010000001;
                8'd042: out <= 14'b11000010000111;
                8'd043: out <= 14'b11000010001110;
                8'd044: out <= 14'b11000010010100;
                8'd045: out <= 14'b11000010011011;
                8'd046: out <= 14'b11000010100010;
                8'd047: out <= 14'b11000010101001;
                8'd048: out <= 14'b11000010110000;
                8'd049: out <= 14'b11000010111000;
                8'd050: out <= 14'b11000010111111;
                8'd051: out <= 14'b11000011000111;
                8'd052: out <= 14'b11000011001111;
                8'd053: out <= 14'b11000011010111;
                8'd054: out <= 14'b11000011011111;
                8'd055: out <= 14'b11000011100111;
                8'd056: out <= 14'b11000011101111;
                8'd057: out <= 14'b11000011111000;
                8'd058: out <= 14'b11000100000001;
                8'd059: out <= 14'b11000100001001;
                8'd060: out <= 14'b11000100010010;
                8'd061: out <= 14'b11000100011100;
                8'd062: out <= 14'b11000100100101;
                8'd063: out <= 14'b11000100101110;
                8'd064: out <= 14'b11000100111000;
                8'd065: out <= 14'b11000101000001;
                8'd066: out <= 14'b11000101001011;
                8'd067: out <= 14'b11000101010101;
                8'd068: out <= 14'b11000101011111;
                8'd069: out <= 14'b11000101101010;
                8'd070: out <= 14'b11000101110100;
                8'd071: out <= 14'b11000101111111;
                8'd072: out <= 14'b11000110001001;
                8'd073: out <= 14'b11000110010100;
                8'd074: out <= 14'b11000110011111;
                8'd075: out <= 14'b11000110101010;
                8'd076: out <= 14'b11000110110101;
                8'd077: out <= 14'b11000111000001;
                8'd078: out <= 14'b11000111001100;
                8'd079: out <= 14'b11000111011000;
                8'd080: out <= 14'b11000111100100;
                8'd081: out <= 14'b11000111110000;
                8'd082: out <= 14'b11000111111100;
                8'd083: out <= 14'b11001000001000;
                8'd084: out <= 14'b11001000010100;
                8'd085: out <= 14'b11001000100001;
                8'd086: out <= 14'b11001000101101;
                8'd087: out <= 14'b11001000111010;
                8'd088: out <= 14'b11001001000111;
                8'd089: out <= 14'b11001001010100;
                8'd090: out <= 14'b11001001100001;
                8'd091: out <= 14'b11001001101110;
                8'd092: out <= 14'b11001001111011;
                8'd093: out <= 14'b11001010001001;
                8'd094: out <= 14'b11001010010111;
                8'd095: out <= 14'b11001010100100;
                8'd096: out <= 14'b11001010110010;
                8'd097: out <= 14'b11001011000000;
                8'd098: out <= 14'b11001011001110;
                8'd099: out <= 14'b11001011011101;
                8'd100: out <= 14'b11001011101011;
                8'd101: out <= 14'b11001011111010;
                8'd102: out <= 14'b11001100001000;
                8'd103: out <= 14'b11001100010111;
                8'd104: out <= 14'b11001100100110;
                8'd105: out <= 14'b11001100110101;
                8'd106: out <= 14'b11001101000100;
                8'd107: out <= 14'b11001101010100;
                8'd108: out <= 14'b11001101100011;
                8'd109: out <= 14'b11001101110010;
                8'd110: out <= 14'b11001110000010;
                8'd111: out <= 14'b11001110010010;
                8'd112: out <= 14'b11001110100010;
                8'd113: out <= 14'b11001110110010;
                8'd114: out <= 14'b11001111000010;
                8'd115: out <= 14'b11001111010010;
                8'd116: out <= 14'b11001111100010;
                8'd117: out <= 14'b11001111110011;
                8'd118: out <= 14'b11010000000100;
                8'd119: out <= 14'b11010000010100;
                8'd120: out <= 14'b11010000100101;
                8'd121: out <= 14'b11010000110110;
                8'd122: out <= 14'b11010001000111;
                8'd123: out <= 14'b11010001011000;
                8'd124: out <= 14'b11010001101001;
                8'd125: out <= 14'b11010001111011;
                8'd126: out <= 14'b11010010001100;
                8'd127: out <= 14'b11010010011110;
                8'd128: out <= 14'b11010010110000;
                8'd129: out <= 14'b11010011000010;
                8'd130: out <= 14'b11010011010011;
                8'd131: out <= 14'b11010011100101;
                8'd132: out <= 14'b11010011111000;
                8'd133: out <= 14'b11010100001010;
                8'd134: out <= 14'b11010100011100;
                8'd135: out <= 14'b11010100101111;
                8'd136: out <= 14'b11010101000001;
                8'd137: out <= 14'b11010101010100;
                8'd138: out <= 14'b11010101100111;
                8'd139: out <= 14'b11010101111010;
                8'd140: out <= 14'b11010110001101;
                8'd141: out <= 14'b11010110100000;
                8'd142: out <= 14'b11010110110011;
                8'd143: out <= 14'b11010111000110;
                8'd144: out <= 14'b11010111011010;
                8'd145: out <= 14'b11010111101101;
                8'd146: out <= 14'b11011000000001;
                8'd147: out <= 14'b11011000010100;
                8'd148: out <= 14'b11011000101000;
                8'd149: out <= 14'b11011000111100;
                8'd150: out <= 14'b11011001010000;
                8'd151: out <= 14'b11011001100100;
                8'd152: out <= 14'b11011001111000;
                8'd153: out <= 14'b11011010001100;
                8'd154: out <= 14'b11011010100001;
                8'd155: out <= 14'b11011010110101;
                8'd156: out <= 14'b11011011001001;
                8'd157: out <= 14'b11011011011110;
                8'd158: out <= 14'b11011011110011;
                8'd159: out <= 14'b11011100001000;
                8'd160: out <= 14'b11011100011100;
                8'd161: out <= 14'b11011100110001;
                8'd162: out <= 14'b11011101000110;
                8'd163: out <= 14'b11011101011011;
                8'd164: out <= 14'b11011101110001;
                8'd165: out <= 14'b11011110000110;
                8'd166: out <= 14'b11011110011011;
                8'd167: out <= 14'b11011110110001;
                8'd168: out <= 14'b11011111000110;
                8'd169: out <= 14'b11011111011100;
                8'd170: out <= 14'b11011111110010;
                8'd171: out <= 14'b11100000000111;
                8'd172: out <= 14'b11100000011101;
                8'd173: out <= 14'b11100000110011;
                8'd174: out <= 14'b11100001001001;
                8'd175: out <= 14'b11100001011111;
                8'd176: out <= 14'b11100001110101;
                8'd177: out <= 14'b11100010001011;
                8'd178: out <= 14'b11100010100010;
                8'd179: out <= 14'b11100010111000;
                8'd180: out <= 14'b11100011001110;
                8'd181: out <= 14'b11100011100101;
                8'd182: out <= 14'b11100011111011;
                8'd183: out <= 14'b11100100010010;
                8'd184: out <= 14'b11100100101001;
                8'd185: out <= 14'b11100100111111;
                8'd186: out <= 14'b11100101010110;
                8'd187: out <= 14'b11100101101101;
                8'd188: out <= 14'b11100110000100;
                8'd189: out <= 14'b11100110011011;
                8'd190: out <= 14'b11100110110010;
                8'd191: out <= 14'b11100111001001;
                8'd192: out <= 14'b11100111100001;
                8'd193: out <= 14'b11100111111000;
                8'd194: out <= 14'b11101000001111;
                8'd195: out <= 14'b11101000100110;
                8'd196: out <= 14'b11101000111110;
                8'd197: out <= 14'b11101001010101;
                8'd198: out <= 14'b11101001101101;
                8'd199: out <= 14'b11101010000100;
                8'd200: out <= 14'b11101010011100;
                8'd201: out <= 14'b11101010110100;
                8'd202: out <= 14'b11101011001100;
                8'd203: out <= 14'b11101011100011;
                8'd204: out <= 14'b11101011111011;
                8'd205: out <= 14'b11101100010011;
                8'd206: out <= 14'b11101100101011;
                8'd207: out <= 14'b11101101000011;
                8'd208: out <= 14'b11101101011011;
                8'd209: out <= 14'b11101101110011;
                8'd210: out <= 14'b11101110001011;
                8'd211: out <= 14'b11101110100011;
                8'd212: out <= 14'b11101110111100;
                8'd213: out <= 14'b11101111010100;
                8'd214: out <= 14'b11101111101100;
                8'd215: out <= 14'b11110000000100;
                8'd216: out <= 14'b11110000011101;
                8'd217: out <= 14'b11110000110101;
                8'd218: out <= 14'b11110001001110;
                8'd219: out <= 14'b11110001100110;
                8'd220: out <= 14'b11110001111111;
                8'd221: out <= 14'b11110010010111;
                8'd222: out <= 14'b11110010110000;
                8'd223: out <= 14'b11110011001000;
                8'd224: out <= 14'b11110011100001;
                8'd225: out <= 14'b11110011111010;
                8'd226: out <= 14'b11110100010010;
                8'd227: out <= 14'b11110100101011;
                8'd228: out <= 14'b11110101000100;
                8'd229: out <= 14'b11110101011101;
                8'd230: out <= 14'b11110101110101;
                8'd231: out <= 14'b11110110001110;
                8'd232: out <= 14'b11110110100111;
                8'd233: out <= 14'b11110111000000;
                8'd234: out <= 14'b11110111011001;
                8'd235: out <= 14'b11110111110010;
                8'd236: out <= 14'b11111000001011;
                8'd237: out <= 14'b11111000100100;
                8'd238: out <= 14'b11111000111101;
                8'd239: out <= 14'b11111001010110;
                8'd240: out <= 14'b11111001101111;
                8'd241: out <= 14'b11111010001000;
                8'd242: out <= 14'b11111010100001;
                8'd243: out <= 14'b11111010111010;
                8'd244: out <= 14'b11111011010011;
                8'd245: out <= 14'b11111011101100;
                8'd246: out <= 14'b11111100000101;
                8'd247: out <= 14'b11111100011110;
                8'd248: out <= 14'b11111100110111;
                8'd249: out <= 14'b11111101010000;
                8'd250: out <= 14'b11111101101001;
                8'd251: out <= 14'b11111110000010;
                8'd252: out <= 14'b11111110011011;
                8'd253: out <= 14'b11111110110101;
                8'd254: out <= 14'b11111111001110;
                8'd255: out <= 14'b11111111100111;
            endcase        end
    endcase
end

endmodule