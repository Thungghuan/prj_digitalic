
module s2p32bit(   //为了后续步骤方便，直接替换原来的移位寄存器工程文件
    input        clk  ,  //系统时钟, 500MHz
 input         [15:0]        a, //整个函数的输入变量
 input [15:0]         b,
 input [4:0]  c,
    output  reg [10:0]  y  //有10位正弦信号的输出, 此时y变为有符号数，最高位为符号位
    );
 
 wire  [9:0]  x; //abc的后10位
 
//wire [21:0] abc; //正弦函数的输入变量（a+b）×c, 一共22位
//reg [5:0] n; //用于排查问题
//assign abc = (a+b)*c; //此处如果一步到位，综合出来的是组合逻辑
 
//以下使用流水线实现乘法器
wire  [16:0] mul_a;  //a和b相加有17位
wire  [4:0] mul_b;   //c只有5位
 reg  [21:0] mul_out; //乘法器的输出, 22位
 
 assign mul_a = a+b;
 assign mul_b = c;
 
reg [21:0] store0,store1,store2,store3,store4;  //用于暂存部分积
reg [21:0] add01, add12, add23;

//将部分积暂存，之后再加
always @ (posedge clk)  begin
store0 <= mul_b[0] ? {5'b0,mul_a}:22'b0;      
 end
 
always @ (posedge clk)  begin
 store1 <= mul_b[1] ? {4'b0,mul_a,1'b0}:22'b0;
add01  <= store1+store0;
 end 

always @ (posedge clk)  begin
 store2 <= mul_b[2] ? {3'b0,mul_a,2'b0}:22'b0;
add12  <= add01+store2;
 end 

always @ (posedge clk)  begin
 store3 <= mul_b[3] ? {2'b0,mul_a,3'b0}:22'b0;
add23  <= add12+store3;
 end 

always @ (posedge clk)  begin
 store4 <= mul_b[3] ? {1'b0,mul_a,4'b0}:22'b0;
mul_out  <= add23+store4;
 end 
 
assign x = mul_out [9:0] ;  
//将乘法结果mul_out的后10位取出来，进入正弦运算，前面的12位不会影响正弦运算的结果
                                                                                                                                                                                                                      
 
always @(posedge clk)  begin   
//此处不再使用ip核或mif文件，直接用case语句查表

case (x)   //三角函数表的深度为1024行，精度为10位
       
		10'd0: y<= 11'b00000000000;
		10'd1: y<= 11'b00000000110;
		10'd2: y<= 11'b00000001101;
		10'd3: y<= 11'b00000010011;
		10'd4: y<= 11'b00000011001;
		10'd5: y<= 11'b00000011111;
		10'd6: y<= 11'b00000100110;
		10'd7: y<= 11'b00000101100;
		10'd8: y<= 11'b00000110010;
		10'd9: y<= 11'b00000111001;
		10'd10: y<= 11'b00000111111;
		10'd11: y<= 11'b00001000101;
		10'd12: y<= 11'b00001001011;
		10'd13: y<= 11'b00001010010;
		10'd14: y<= 11'b00001011000;
		10'd15: y<= 11'b00001011110;
		10'd16: y<= 11'b00001100100;
		10'd17: y<= 11'b00001101011;
		10'd18: y<= 11'b00001110001;
		10'd19: y<= 11'b00001110111;
		10'd20: y<= 11'b00001111101;
		10'd21: y<= 11'b00010000100;
		10'd22: y<= 11'b00010001010;
		10'd23: y<= 11'b00010010000;
		10'd24: y<= 11'b00010010110;
		10'd25: y<= 11'b00010011100;
		10'd26: y<= 11'b00010100011;
		10'd27: y<= 11'b00010101001;
		10'd28: y<= 11'b00010101111;
		10'd29: y<= 11'b00010110101;
		10'd30: y<= 11'b00010111011;
		10'd31: y<= 11'b00011000010;
		10'd32: y<= 11'b00011001000;
		10'd33: y<= 11'b00011001110;
		10'd34: y<= 11'b00011010100;
		10'd35: y<= 11'b00011011010;
		10'd36: y<= 11'b00011100000;
		10'd37: y<= 11'b00011100110;
		10'd38: y<= 11'b00011101101;
		10'd39: y<= 11'b00011110011;
		10'd40: y<= 11'b00011111001;
		10'd41: y<= 11'b00011111111;
		10'd42: y<= 11'b00100000101;
		10'd43: y<= 11'b00100001011;
		10'd44: y<= 11'b00100010001;
		10'd45: y<= 11'b00100010111;
		10'd46: y<= 11'b00100011101;
		10'd47: y<= 11'b00100100011;
		10'd48: y<= 11'b00100101001;
		10'd49: y<= 11'b00100101111;
		10'd50: y<= 11'b00100110101;
		10'd51: y<= 11'b00100111011;
		10'd52: y<= 11'b00101000001;
		10'd53: y<= 11'b00101000111;
		10'd54: y<= 11'b00101001101;
		10'd55: y<= 11'b00101010011;
		10'd56: y<= 11'b00101011001;
		10'd57: y<= 11'b00101011111;
		10'd58: y<= 11'b00101100101;
		10'd59: y<= 11'b00101101011;
		10'd60: y<= 11'b00101110001;
		10'd61: y<= 11'b00101110110;
		10'd62: y<= 11'b00101111100;
		10'd63: y<= 11'b00110000010;
		10'd64: y<= 11'b00110001000;
		10'd65: y<= 11'b00110001110;
		10'd66: y<= 11'b00110010011;
		10'd67: y<= 11'b00110011001;
		10'd68: y<= 11'b00110011111;
		10'd69: y<= 11'b00110100101;
		10'd70: y<= 11'b00110101010;
		10'd71: y<= 11'b00110110000;
		10'd72: y<= 11'b00110110110;
		10'd73: y<= 11'b00110111011;
		10'd74: y<= 11'b00111000001;
		10'd75: y<= 11'b00111000111;
		10'd76: y<= 11'b00111001100;
		10'd77: y<= 11'b00111010010;
		10'd78: y<= 11'b00111011000;
		10'd79: y<= 11'b00111011101;
		10'd80: y<= 11'b00111100011;
		10'd81: y<= 11'b00111101000;
		10'd82: y<= 11'b00111101110;
		10'd83: y<= 11'b00111110011;
		10'd84: y<= 11'b00111111001;
		10'd85: y<= 11'b00111111110;
		10'd86: y<= 11'b01000000100;
		10'd87: y<= 11'b01000001001;
		10'd88: y<= 11'b01000001110;
		10'd89: y<= 11'b01000010100;
		10'd90: y<= 11'b01000011001;
		10'd91: y<= 11'b01000011111;
		10'd92: y<= 11'b01000100100;
		10'd93: y<= 11'b01000101001;
		10'd94: y<= 11'b01000101110;
		10'd95: y<= 11'b01000110100;
		10'd96: y<= 11'b01000111001;
		10'd97: y<= 11'b01000111110;
		10'd98: y<= 11'b01001000011;
		10'd99: y<= 11'b01001001000;
		10'd100: y<= 11'b01001001110;
		10'd101: y<= 11'b01001010011;
		10'd102: y<= 11'b01001011000;
		10'd103: y<= 11'b01001011101;
		10'd104: y<= 11'b01001100010;
		10'd105: y<= 11'b01001100111;
		10'd106: y<= 11'b01001101100;
		10'd107: y<= 11'b01001110001;
		10'd108: y<= 11'b01001110110;
		10'd109: y<= 11'b01001111011;
		10'd110: y<= 11'b01010000000;
		10'd111: y<= 11'b01010000101;
		10'd112: y<= 11'b01010001010;
		10'd113: y<= 11'b01010001110;
		10'd114: y<= 11'b01010010011;
		10'd115: y<= 11'b01010011000;
		10'd116: y<= 11'b01010011101;
		10'd117: y<= 11'b01010100010;
		10'd118: y<= 11'b01010100110;
		10'd119: y<= 11'b01010101011;
		10'd120: y<= 11'b01010110000;
		10'd121: y<= 11'b01010110100;
		10'd122: y<= 11'b01010111001;
		10'd123: y<= 11'b01010111110;
		10'd124: y<= 11'b01011000010;
		10'd125: y<= 11'b01011000111;
		10'd126: y<= 11'b01011001011;
		10'd127: y<= 11'b01011010000;
		10'd128: y<= 11'b01011010100;
		10'd129: y<= 11'b01011011001;
		10'd130: y<= 11'b01011011101;
		10'd131: y<= 11'b01011100001;
		10'd132: y<= 11'b01011100110;
		10'd133: y<= 11'b01011101010;
		10'd134: y<= 11'b01011101110;
		10'd135: y<= 11'b01011110011;
		10'd136: y<= 11'b01011110111;
		10'd137: y<= 11'b01011111011;
		10'd138: y<= 11'b01011111111;
		10'd139: y<= 11'b01100000011;
		10'd140: y<= 11'b01100000111;
		10'd141: y<= 11'b01100001011;
		10'd142: y<= 11'b01100010000;
		10'd143: y<= 11'b01100010100;
		10'd144: y<= 11'b01100011000;
		10'd145: y<= 11'b01100011100;
		10'd146: y<= 11'b01100011111;
		10'd147: y<= 11'b01100100011;
		10'd148: y<= 11'b01100100111;
		10'd149: y<= 11'b01100101011;
		10'd150: y<= 11'b01100101111;
		10'd151: y<= 11'b01100110011;
		10'd152: y<= 11'b01100110110;
		10'd153: y<= 11'b01100111010;
		10'd154: y<= 11'b01100111110;
		10'd155: y<= 11'b01101000010;
		10'd156: y<= 11'b01101000101;
		10'd157: y<= 11'b01101001001;
		10'd158: y<= 11'b01101001100;
		10'd159: y<= 11'b01101010000;
		10'd160: y<= 11'b01101010011;
		10'd161: y<= 11'b01101010111;
		10'd162: y<= 11'b01101011010;
		10'd163: y<= 11'b01101011110;
		10'd164: y<= 11'b01101100001;
		10'd165: y<= 11'b01101100100;
		10'd166: y<= 11'b01101101000;
		10'd167: y<= 11'b01101101011;
		10'd168: y<= 11'b01101101110;
		10'd169: y<= 11'b01101110010;
		10'd170: y<= 11'b01101110101;
		10'd171: y<= 11'b01101111000;
		10'd172: y<= 11'b01101111011;
		10'd173: y<= 11'b01101111110;
		10'd174: y<= 11'b01110000001;
		10'd175: y<= 11'b01110000100;
		10'd176: y<= 11'b01110000111;
		10'd177: y<= 11'b01110001010;
		10'd178: y<= 11'b01110001101;
		10'd179: y<= 11'b01110010000;
		10'd180: y<= 11'b01110010011;
		10'd181: y<= 11'b01110010101;
		10'd182: y<= 11'b01110011000;
		10'd183: y<= 11'b01110011011;
		10'd184: y<= 11'b01110011110;
		10'd185: y<= 11'b01110100000;
		10'd186: y<= 11'b01110100011;
		10'd187: y<= 11'b01110100110;
		10'd188: y<= 11'b01110101000;
		10'd189: y<= 11'b01110101011;
		10'd190: y<= 11'b01110101101;
		10'd191: y<= 11'b01110110000;
		10'd192: y<= 11'b01110110010;
		10'd193: y<= 11'b01110110100;
		10'd194: y<= 11'b01110110111;
		10'd195: y<= 11'b01110111001;
		10'd196: y<= 11'b01110111011;
		10'd197: y<= 11'b01110111110;
		10'd198: y<= 11'b01111000000;
		10'd199: y<= 11'b01111000010;
		10'd200: y<= 11'b01111000100;
		10'd201: y<= 11'b01111000110;
		10'd202: y<= 11'b01111001000;
		10'd203: y<= 11'b01111001010;
		10'd204: y<= 11'b01111001100;
		10'd205: y<= 11'b01111001110;
		10'd206: y<= 11'b01111010000;
		10'd207: y<= 11'b01111010010;
		10'd208: y<= 11'b01111010100;
		10'd209: y<= 11'b01111010110;
		10'd210: y<= 11'b01111010111;
		10'd211: y<= 11'b01111011001;
		10'd212: y<= 11'b01111011011;
		10'd213: y<= 11'b01111011101;
		10'd214: y<= 11'b01111011110;
		10'd215: y<= 11'b01111100000;
		10'd216: y<= 11'b01111100001;
		10'd217: y<= 11'b01111100011;
		10'd218: y<= 11'b01111100100;
		10'd219: y<= 11'b01111100110;
		10'd220: y<= 11'b01111100111;
		10'd221: y<= 11'b01111101000;
		10'd222: y<= 11'b01111101010;
		10'd223: y<= 11'b01111101011;
		10'd224: y<= 11'b01111101100;
		10'd225: y<= 11'b01111101110;
		10'd226: y<= 11'b01111101111;
		10'd227: y<= 11'b01111110000;
		10'd228: y<= 11'b01111110001;
		10'd229: y<= 11'b01111110010;
		10'd230: y<= 11'b01111110011;
		10'd231: y<= 11'b01111110100;
		10'd232: y<= 11'b01111110101;
		10'd233: y<= 11'b01111110110;
		10'd234: y<= 11'b01111110111;
		10'd235: y<= 11'b01111111000;
		10'd236: y<= 11'b01111111000;
		10'd237: y<= 11'b01111111001;
		10'd238: y<= 11'b01111111010;
		10'd239: y<= 11'b01111111010;
		10'd240: y<= 11'b01111111011;
		10'd241: y<= 11'b01111111100;
		10'd242: y<= 11'b01111111100;
		10'd243: y<= 11'b01111111101;
		10'd244: y<= 11'b01111111101;
		10'd245: y<= 11'b01111111110;
		10'd246: y<= 11'b01111111110;
		10'd247: y<= 11'b01111111110;
		10'd248: y<= 11'b01111111111;
		10'd249: y<= 11'b01111111111;
		10'd250: y<= 11'b01111111111;
		10'd251: y<= 11'b01111111111;
		10'd252: y<= 11'b01111111111;
		10'd253: y<= 11'b01111111111;
		10'd254: y<= 11'b01111111111;
		10'd255: y<= 11'b01111111111;
		10'd256: y<= 11'b01111111111;
		10'd257: y<= 11'b01111111111;
		10'd258: y<= 11'b01111111111;
		10'd259: y<= 11'b01111111111;
		10'd260: y<= 11'b01111111111;
		10'd261: y<= 11'b01111111111;
		10'd262: y<= 11'b01111111111;
		10'd263: y<= 11'b01111111111;
		10'd264: y<= 11'b01111111111;
		10'd265: y<= 11'b01111111110;
		10'd266: y<= 11'b01111111110;
		10'd267: y<= 11'b01111111110;
		10'd268: y<= 11'b01111111101;
		10'd269: y<= 11'b01111111101;
		10'd270: y<= 11'b01111111100;
		10'd271: y<= 11'b01111111100;
		10'd272: y<= 11'b01111111011;
		10'd273: y<= 11'b01111111010;
		10'd274: y<= 11'b01111111010;
		10'd275: y<= 11'b01111111001;
		10'd276: y<= 11'b01111111000;
		10'd277: y<= 11'b01111111000;
		10'd278: y<= 11'b01111110111;
		10'd279: y<= 11'b01111110110;
		10'd280: y<= 11'b01111110101;
		10'd281: y<= 11'b01111110100;
		10'd282: y<= 11'b01111110011;
		10'd283: y<= 11'b01111110010;
		10'd284: y<= 11'b01111110001;
		10'd285: y<= 11'b01111110000;
		10'd286: y<= 11'b01111101111;
		10'd287: y<= 11'b01111101110;
		10'd288: y<= 11'b01111101100;
		10'd289: y<= 11'b01111101011;
		10'd290: y<= 11'b01111101010;
		10'd291: y<= 11'b01111101000;
		10'd292: y<= 11'b01111100111;
		10'd293: y<= 11'b01111100110;
		10'd294: y<= 11'b01111100100;
		10'd295: y<= 11'b01111100011;
		10'd296: y<= 11'b01111100001;
		10'd297: y<= 11'b01111100000;
		10'd298: y<= 11'b01111011110;
		10'd299: y<= 11'b01111011101;
		10'd300: y<= 11'b01111011011;
		10'd301: y<= 11'b01111011001;
		10'd302: y<= 11'b01111010111;
		10'd303: y<= 11'b01111010110;
		10'd304: y<= 11'b01111010100;
		10'd305: y<= 11'b01111010010;
		10'd306: y<= 11'b01111010000;
		10'd307: y<= 11'b01111001110;
		10'd308: y<= 11'b01111001100;
		10'd309: y<= 11'b01111001010;
		10'd310: y<= 11'b01111001000;
		10'd311: y<= 11'b01111000110;
		10'd312: y<= 11'b01111000100;
		10'd313: y<= 11'b01111000010;
		10'd314: y<= 11'b01111000000;
		10'd315: y<= 11'b01110111110;
		10'd316: y<= 11'b01110111011;
		10'd317: y<= 11'b01110111001;
		10'd318: y<= 11'b01110110111;
		10'd319: y<= 11'b01110110100;
		10'd320: y<= 11'b01110110010;
		10'd321: y<= 11'b01110110000;
		10'd322: y<= 11'b01110101101;
		10'd323: y<= 11'b01110101011;
		10'd324: y<= 11'b01110101000;
		10'd325: y<= 11'b01110100110;
		10'd326: y<= 11'b01110100011;
		10'd327: y<= 11'b01110100000;
		10'd328: y<= 11'b01110011110;
		10'd329: y<= 11'b01110011011;
		10'd330: y<= 11'b01110011000;
		10'd331: y<= 11'b01110010101;
		10'd332: y<= 11'b01110010011;
		10'd333: y<= 11'b01110010000;
		10'd334: y<= 11'b01110001101;
		10'd335: y<= 11'b01110001010;
		10'd336: y<= 11'b01110000111;
		10'd337: y<= 11'b01110000100;
		10'd338: y<= 11'b01110000001;
		10'd339: y<= 11'b01101111110;
		10'd340: y<= 11'b01101111011;
		10'd341: y<= 11'b01101111000;
		10'd342: y<= 11'b01101110101;
		10'd343: y<= 11'b01101110010;
		10'd344: y<= 11'b01101101110;
		10'd345: y<= 11'b01101101011;
		10'd346: y<= 11'b01101101000;
		10'd347: y<= 11'b01101100100;
		10'd348: y<= 11'b01101100001;
		10'd349: y<= 11'b01101011110;
		10'd350: y<= 11'b01101011010;
		10'd351: y<= 11'b01101010111;
		10'd352: y<= 11'b01101010011;
		10'd353: y<= 11'b01101010000;
		10'd354: y<= 11'b01101001100;
		10'd355: y<= 11'b01101001001;
		10'd356: y<= 11'b01101000101;
		10'd357: y<= 11'b01101000010;
		10'd358: y<= 11'b01100111110;
		10'd359: y<= 11'b01100111010;
		10'd360: y<= 11'b01100110110;
		10'd361: y<= 11'b01100110011;
		10'd362: y<= 11'b01100101111;
		10'd363: y<= 11'b01100101011;
		10'd364: y<= 11'b01100100111;
		10'd365: y<= 11'b01100100011;
		10'd366: y<= 11'b01100011111;
		10'd367: y<= 11'b01100011100;
		10'd368: y<= 11'b01100011000;
		10'd369: y<= 11'b01100010100;
		10'd370: y<= 11'b01100010000;
		10'd371: y<= 11'b01100001011;
		10'd372: y<= 11'b01100000111;
		10'd373: y<= 11'b01100000011;
		10'd374: y<= 11'b01011111111;
		10'd375: y<= 11'b01011111011;
		10'd376: y<= 11'b01011110111;
		10'd377: y<= 11'b01011110011;
		10'd378: y<= 11'b01011101110;
		10'd379: y<= 11'b01011101010;
		10'd380: y<= 11'b01011100110;
		10'd381: y<= 11'b01011100001;
		10'd382: y<= 11'b01011011101;
		10'd383: y<= 11'b01011011001;
		10'd384: y<= 11'b01011010100;
		10'd385: y<= 11'b01011010000;
		10'd386: y<= 11'b01011001011;
		10'd387: y<= 11'b01011000111;
		10'd388: y<= 11'b01011000010;
		10'd389: y<= 11'b01010111110;
		10'd390: y<= 11'b01010111001;
		10'd391: y<= 11'b01010110100;
		10'd392: y<= 11'b01010110000;
		10'd393: y<= 11'b01010101011;
		10'd394: y<= 11'b01010100110;
		10'd395: y<= 11'b01010100010;
		10'd396: y<= 11'b01010011101;
		10'd397: y<= 11'b01010011000;
		10'd398: y<= 11'b01010010011;
		10'd399: y<= 11'b01010001110;
		10'd400: y<= 11'b01010001010;
		10'd401: y<= 11'b01010000101;
		10'd402: y<= 11'b01010000000;
		10'd403: y<= 11'b01001111011;
		10'd404: y<= 11'b01001110110;
		10'd405: y<= 11'b01001110001;
		10'd406: y<= 11'b01001101100;
		10'd407: y<= 11'b01001100111;
		10'd408: y<= 11'b01001100010;
		10'd409: y<= 11'b01001011101;
		10'd410: y<= 11'b01001011000;
		10'd411: y<= 11'b01001010011;
		10'd412: y<= 11'b01001001110;
		10'd413: y<= 11'b01001001000;
		10'd414: y<= 11'b01001000011;
		10'd415: y<= 11'b01000111110;
		10'd416: y<= 11'b01000111001;
		10'd417: y<= 11'b01000110100;
		10'd418: y<= 11'b01000101110;
		10'd419: y<= 11'b01000101001;
		10'd420: y<= 11'b01000100100;
		10'd421: y<= 11'b01000011111;
		10'd422: y<= 11'b01000011001;
		10'd423: y<= 11'b01000010100;
		10'd424: y<= 11'b01000001110;
		10'd425: y<= 11'b01000001001;
		10'd426: y<= 11'b01000000100;
		10'd427: y<= 11'b00111111110;
		10'd428: y<= 11'b00111111001;
		10'd429: y<= 11'b00111110011;
		10'd430: y<= 11'b00111101110;
		10'd431: y<= 11'b00111101000;
		10'd432: y<= 11'b00111100011;
		10'd433: y<= 11'b00111011101;
		10'd434: y<= 11'b00111011000;
		10'd435: y<= 11'b00111010010;
		10'd436: y<= 11'b00111001100;
		10'd437: y<= 11'b00111000111;
		10'd438: y<= 11'b00111000001;
		10'd439: y<= 11'b00110111011;
		10'd440: y<= 11'b00110110110;
		10'd441: y<= 11'b00110110000;
		10'd442: y<= 11'b00110101010;
		10'd443: y<= 11'b00110100101;
		10'd444: y<= 11'b00110011111;
		10'd445: y<= 11'b00110011001;
		10'd446: y<= 11'b00110010011;
		10'd447: y<= 11'b00110001110;
		10'd448: y<= 11'b00110001000;
		10'd449: y<= 11'b00110000010;
		10'd450: y<= 11'b00101111100;
		10'd451: y<= 11'b00101110110;
		10'd452: y<= 11'b00101110001;
		10'd453: y<= 11'b00101101011;
		10'd454: y<= 11'b00101100101;
		10'd455: y<= 11'b00101011111;
		10'd456: y<= 11'b00101011001;
		10'd457: y<= 11'b00101010011;
		10'd458: y<= 11'b00101001101;
		10'd459: y<= 11'b00101000111;
		10'd460: y<= 11'b00101000001;
		10'd461: y<= 11'b00100111011;
		10'd462: y<= 11'b00100110101;
		10'd463: y<= 11'b00100101111;
		10'd464: y<= 11'b00100101001;
		10'd465: y<= 11'b00100100011;
		10'd466: y<= 11'b00100011101;
		10'd467: y<= 11'b00100010111;
		10'd468: y<= 11'b00100010001;
		10'd469: y<= 11'b00100001011;
		10'd470: y<= 11'b00100000101;
		10'd471: y<= 11'b00011111111;
		10'd472: y<= 11'b00011111001;
		10'd473: y<= 11'b00011110011;
		10'd474: y<= 11'b00011101101;
		10'd475: y<= 11'b00011100110;
		10'd476: y<= 11'b00011100000;
		10'd477: y<= 11'b00011011010;
		10'd478: y<= 11'b00011010100;
		10'd479: y<= 11'b00011001110;
		10'd480: y<= 11'b00011001000;
		10'd481: y<= 11'b00011000010;
		10'd482: y<= 11'b00010111011;
		10'd483: y<= 11'b00010110101;
		10'd484: y<= 11'b00010101111;
		10'd485: y<= 11'b00010101001;
		10'd486: y<= 11'b00010100011;
		10'd487: y<= 11'b00010011100;
		10'd488: y<= 11'b00010010110;
		10'd489: y<= 11'b00010010000;
		10'd490: y<= 11'b00010001010;
		10'd491: y<= 11'b00010000100;
		10'd492: y<= 11'b00001111101;
		10'd493: y<= 11'b00001110111;
		10'd494: y<= 11'b00001110001;
		10'd495: y<= 11'b00001101011;
		10'd496: y<= 11'b00001100100;
		10'd497: y<= 11'b00001011110;
		10'd498: y<= 11'b00001011000;
		10'd499: y<= 11'b00001010010;
		10'd500: y<= 11'b00001001011;
		10'd501: y<= 11'b00001000101;
		10'd502: y<= 11'b00000111111;
		10'd503: y<= 11'b00000111001;
		10'd504: y<= 11'b00000110010;
		10'd505: y<= 11'b00000101100;
		10'd506: y<= 11'b00000100110;
		10'd507: y<= 11'b00000011111;
		10'd508: y<= 11'b00000011001;
		10'd509: y<= 11'b00000010011;
		10'd510: y<= 11'b00000001101;
		10'd511: y<= 11'b00000000110;
		10'd512: y<= 11'b00000000000;
		10'd513: y<= 11'b11111111010;
		10'd514: y<= 11'b11111110011;
		10'd515: y<= 11'b11111101101;
		10'd516: y<= 11'b11111100111;
		10'd517: y<= 11'b11111100001;
		10'd518: y<= 11'b11111011010;
		10'd519: y<= 11'b11111010100;
		10'd520: y<= 11'b11111001110;
		10'd521: y<= 11'b11111000111;
		10'd522: y<= 11'b11111000001;
		10'd523: y<= 11'b11110111011;
		10'd524: y<= 11'b11110110101;
		10'd525: y<= 11'b11110101110;
		10'd526: y<= 11'b11110101000;
		10'd527: y<= 11'b11110100010;
		10'd528: y<= 11'b11110011100;
		10'd529: y<= 11'b11110010101;
		10'd530: y<= 11'b11110001111;
		10'd531: y<= 11'b11110001001;
		10'd532: y<= 11'b11110000011;
		10'd533: y<= 11'b11101111100;
		10'd534: y<= 11'b11101110110;
		10'd535: y<= 11'b11101110000;
		10'd536: y<= 11'b11101101010;
		10'd537: y<= 11'b11101100100;
		10'd538: y<= 11'b11101011101;
		10'd539: y<= 11'b11101010111;
		10'd540: y<= 11'b11101010001;
		10'd541: y<= 11'b11101001011;
		10'd542: y<= 11'b11101000101;
		10'd543: y<= 11'b11100111110;
		10'd544: y<= 11'b11100111000;
		10'd545: y<= 11'b11100110010;
		10'd546: y<= 11'b11100101100;
		10'd547: y<= 11'b11100100110;
		10'd548: y<= 11'b11100100000;
		10'd549: y<= 11'b11100011010;
		10'd550: y<= 11'b11100010011;
		10'd551: y<= 11'b11100001101;
		10'd552: y<= 11'b11100000111;
		10'd553: y<= 11'b11100000001;
		10'd554: y<= 11'b11011111011;
		10'd555: y<= 11'b11011110101;
		10'd556: y<= 11'b11011101111;
		10'd557: y<= 11'b11011101001;
		10'd558: y<= 11'b11011100011;
		10'd559: y<= 11'b11011011101;
		10'd560: y<= 11'b11011010111;
		10'd561: y<= 11'b11011010001;
		10'd562: y<= 11'b11011001011;
		10'd563: y<= 11'b11011000101;
		10'd564: y<= 11'b11010111111;
		10'd565: y<= 11'b11010111001;
		10'd566: y<= 11'b11010110011;
		10'd567: y<= 11'b11010101101;
		10'd568: y<= 11'b11010100111;
		10'd569: y<= 11'b11010100001;
		10'd570: y<= 11'b11010011011;
		10'd571: y<= 11'b11010010101;
		10'd572: y<= 11'b11010001111;
		10'd573: y<= 11'b11010001010;
		10'd574: y<= 11'b11010000100;
		10'd575: y<= 11'b11001111110;
		10'd576: y<= 11'b11001111000;
		10'd577: y<= 11'b11001110010;
		10'd578: y<= 11'b11001101101;
		10'd579: y<= 11'b11001100111;
		10'd580: y<= 11'b11001100001;
		10'd581: y<= 11'b11001011011;
		10'd582: y<= 11'b11001010110;
		10'd583: y<= 11'b11001010000;
		10'd584: y<= 11'b11001001010;
		10'd585: y<= 11'b11001000101;
		10'd586: y<= 11'b11000111111;
		10'd587: y<= 11'b11000111001;
		10'd588: y<= 11'b11000110100;
		10'd589: y<= 11'b11000101110;
		10'd590: y<= 11'b11000101000;
		10'd591: y<= 11'b11000100011;
		10'd592: y<= 11'b11000011101;
		10'd593: y<= 11'b11000011000;
		10'd594: y<= 11'b11000010010;
		10'd595: y<= 11'b11000001101;
		10'd596: y<= 11'b11000000111;
		10'd597: y<= 11'b11000000010;
		10'd598: y<= 11'b10111111100;
		10'd599: y<= 11'b10111110111;
		10'd600: y<= 11'b10111110010;
		10'd601: y<= 11'b10111101100;
		10'd602: y<= 11'b10111100111;
		10'd603: y<= 11'b10111100001;
		10'd604: y<= 11'b10111011100;
		10'd605: y<= 11'b10111010111;
		10'd606: y<= 11'b10111010010;
		10'd607: y<= 11'b10111001100;
		10'd608: y<= 11'b10111000111;
		10'd609: y<= 11'b10111000010;
		10'd610: y<= 11'b10110111101;
		10'd611: y<= 11'b10110111000;
		10'd612: y<= 11'b10110110010;
		10'd613: y<= 11'b10110101101;
		10'd614: y<= 11'b10110101000;
		10'd615: y<= 11'b10110100011;
		10'd616: y<= 11'b10110011110;
		10'd617: y<= 11'b10110011001;
		10'd618: y<= 11'b10110010100;
		10'd619: y<= 11'b10110001111;
		10'd620: y<= 11'b10110001010;
		10'd621: y<= 11'b10110000101;
		10'd622: y<= 11'b10110000000;
		10'd623: y<= 11'b10101111011;
		10'd624: y<= 11'b10101110110;
		10'd625: y<= 11'b10101110010;
		10'd626: y<= 11'b10101101101;
		10'd627: y<= 11'b10101101000;
		10'd628: y<= 11'b10101100011;
		10'd629: y<= 11'b10101011110;
		10'd630: y<= 11'b10101011010;
		10'd631: y<= 11'b10101010101;
		10'd632: y<= 11'b10101010000;
		10'd633: y<= 11'b10101001100;
		10'd634: y<= 11'b10101000111;
		10'd635: y<= 11'b10101000010;
		10'd636: y<= 11'b10100111110;
		10'd637: y<= 11'b10100111001;
		10'd638: y<= 11'b10100110101;
		10'd639: y<= 11'b10100110000;
		10'd640: y<= 11'b10100101100;
		10'd641: y<= 11'b10100100111;
		10'd642: y<= 11'b10100100011;
		10'd643: y<= 11'b10100011111;
		10'd644: y<= 11'b10100011010;
		10'd645: y<= 11'b10100010110;
		10'd646: y<= 11'b10100010010;
		10'd647: y<= 11'b10100001101;
		10'd648: y<= 11'b10100001001;
		10'd649: y<= 11'b10100000101;
		10'd650: y<= 11'b10100000001;
		10'd651: y<= 11'b10011111101;
		10'd652: y<= 11'b10011111001;
		10'd653: y<= 11'b10011110101;
		10'd654: y<= 11'b10011110000;
		10'd655: y<= 11'b10011101100;
		10'd656: y<= 11'b10011101000;
		10'd657: y<= 11'b10011100100;
		10'd658: y<= 11'b10011100001;
		10'd659: y<= 11'b10011011101;
		10'd660: y<= 11'b10011011001;
		10'd661: y<= 11'b10011010101;
		10'd662: y<= 11'b10011010001;
		10'd663: y<= 11'b10011001101;
		10'd664: y<= 11'b10011001010;
		10'd665: y<= 11'b10011000110;
		10'd666: y<= 11'b10011000010;
		10'd667: y<= 11'b10010111110;
		10'd668: y<= 11'b10010111011;
		10'd669: y<= 11'b10010110111;
		10'd670: y<= 11'b10010110100;
		10'd671: y<= 11'b10010110000;
		10'd672: y<= 11'b10010101101;
		10'd673: y<= 11'b10010101001;
		10'd674: y<= 11'b10010100110;
		10'd675: y<= 11'b10010100010;
		10'd676: y<= 11'b10010011111;
		10'd677: y<= 11'b10010011100;
		10'd678: y<= 11'b10010011000;
		10'd679: y<= 11'b10010010101;
		10'd680: y<= 11'b10010010010;
		10'd681: y<= 11'b10010001110;
		10'd682: y<= 11'b10010001011;
		10'd683: y<= 11'b10010001000;
		10'd684: y<= 11'b10010000101;
		10'd685: y<= 11'b10010000010;
		10'd686: y<= 11'b10001111111;
		10'd687: y<= 11'b10001111100;
		10'd688: y<= 11'b10001111001;
		10'd689: y<= 11'b10001110110;
		10'd690: y<= 11'b10001110011;
		10'd691: y<= 11'b10001110000;
		10'd692: y<= 11'b10001101101;
		10'd693: y<= 11'b10001101011;
		10'd694: y<= 11'b10001101000;
		10'd695: y<= 11'b10001100101;
		10'd696: y<= 11'b10001100010;
		10'd697: y<= 11'b10001100000;
		10'd698: y<= 11'b10001011101;
		10'd699: y<= 11'b10001011010;
		10'd700: y<= 11'b10001011000;
		10'd701: y<= 11'b10001010101;
		10'd702: y<= 11'b10001010011;
		10'd703: y<= 11'b10001010000;
		10'd704: y<= 11'b10001001110;
		10'd705: y<= 11'b10001001100;
		10'd706: y<= 11'b10001001001;
		10'd707: y<= 11'b10001000111;
		10'd708: y<= 11'b10001000101;
		10'd709: y<= 11'b10001000010;
		10'd710: y<= 11'b10001000000;
		10'd711: y<= 11'b10000111110;
		10'd712: y<= 11'b10000111100;
		10'd713: y<= 11'b10000111010;
		10'd714: y<= 11'b10000111000;
		10'd715: y<= 11'b10000110110;
		10'd716: y<= 11'b10000110100;
		10'd717: y<= 11'b10000110010;
		10'd718: y<= 11'b10000110000;
		10'd719: y<= 11'b10000101110;
		10'd720: y<= 11'b10000101100;
		10'd721: y<= 11'b10000101010;
		10'd722: y<= 11'b10000101001;
		10'd723: y<= 11'b10000100111;
		10'd724: y<= 11'b10000100101;
		10'd725: y<= 11'b10000100011;
		10'd726: y<= 11'b10000100010;
		10'd727: y<= 11'b10000100000;
		10'd728: y<= 11'b10000011111;
		10'd729: y<= 11'b10000011101;
		10'd730: y<= 11'b10000011100;
		10'd731: y<= 11'b10000011010;
		10'd732: y<= 11'b10000011001;
		10'd733: y<= 11'b10000011000;
		10'd734: y<= 11'b10000010110;
		10'd735: y<= 11'b10000010101;
		10'd736: y<= 11'b10000010100;
		10'd737: y<= 11'b10000010010;
		10'd738: y<= 11'b10000010001;
		10'd739: y<= 11'b10000010000;
		10'd740: y<= 11'b10000001111;
		10'd741: y<= 11'b10000001110;
		10'd742: y<= 11'b10000001101;
		10'd743: y<= 11'b10000001100;
		10'd744: y<= 11'b10000001011;
		10'd745: y<= 11'b10000001010;
		10'd746: y<= 11'b10000001001;
		10'd747: y<= 11'b10000001000;
		10'd748: y<= 11'b10000001000;
		10'd749: y<= 11'b10000000111;
		10'd750: y<= 11'b10000000110;
		10'd751: y<= 11'b10000000110;
		10'd752: y<= 11'b10000000101;
		10'd753: y<= 11'b10000000100;
		10'd754: y<= 11'b10000000100;
		10'd755: y<= 11'b10000000011;
		10'd756: y<= 11'b10000000011;
		10'd757: y<= 11'b10000000010;
		10'd758: y<= 11'b10000000010;
		10'd759: y<= 11'b10000000010;
		10'd760: y<= 11'b10000000001;
		10'd761: y<= 11'b10000000001;
		10'd762: y<= 11'b10000000001;
		10'd763: y<= 11'b10000000000;
		10'd764: y<= 11'b10000000000;
		10'd765: y<= 11'b10000000000;
		10'd766: y<= 11'b10000000000;
		10'd767: y<= 11'b10000000000;
		10'd768: y<= 11'b10000000000;
		10'd769: y<= 11'b10000000000;
		10'd770: y<= 11'b10000000000;
		10'd771: y<= 11'b10000000000;
		10'd772: y<= 11'b10000000000;
		10'd773: y<= 11'b10000000000;
		10'd774: y<= 11'b10000000001;
		10'd775: y<= 11'b10000000001;
		10'd776: y<= 11'b10000000001;
		10'd777: y<= 11'b10000000010;
		10'd778: y<= 11'b10000000010;
		10'd779: y<= 11'b10000000010;
		10'd780: y<= 11'b10000000011;
		10'd781: y<= 11'b10000000011;
		10'd782: y<= 11'b10000000100;
		10'd783: y<= 11'b10000000100;
		10'd784: y<= 11'b10000000101;
		10'd785: y<= 11'b10000000110;
		10'd786: y<= 11'b10000000110;
		10'd787: y<= 11'b10000000111;
		10'd788: y<= 11'b10000001000;
		10'd789: y<= 11'b10000001000;
		10'd790: y<= 11'b10000001001;
		10'd791: y<= 11'b10000001010;
		10'd792: y<= 11'b10000001011;
		10'd793: y<= 11'b10000001100;
		10'd794: y<= 11'b10000001101;
		10'd795: y<= 11'b10000001110;
		10'd796: y<= 11'b10000001111;
		10'd797: y<= 11'b10000010000;
		10'd798: y<= 11'b10000010001;
		10'd799: y<= 11'b10000010010;
		10'd800: y<= 11'b10000010100;
		10'd801: y<= 11'b10000010101;
		10'd802: y<= 11'b10000010110;
		10'd803: y<= 11'b10000011000;
		10'd804: y<= 11'b10000011001;
		10'd805: y<= 11'b10000011010;
		10'd806: y<= 11'b10000011100;
		10'd807: y<= 11'b10000011101;
		10'd808: y<= 11'b10000011111;
		10'd809: y<= 11'b10000100000;
		10'd810: y<= 11'b10000100010;
		10'd811: y<= 11'b10000100011;
		10'd812: y<= 11'b10000100101;
		10'd813: y<= 11'b10000100111;
		10'd814: y<= 11'b10000101001;
		10'd815: y<= 11'b10000101010;
		10'd816: y<= 11'b10000101100;
		10'd817: y<= 11'b10000101110;
		10'd818: y<= 11'b10000110000;
		10'd819: y<= 11'b10000110010;
		10'd820: y<= 11'b10000110100;
		10'd821: y<= 11'b10000110110;
		10'd822: y<= 11'b10000111000;
		10'd823: y<= 11'b10000111010;
		10'd824: y<= 11'b10000111100;
		10'd825: y<= 11'b10000111110;
		10'd826: y<= 11'b10001000000;
		10'd827: y<= 11'b10001000010;
		10'd828: y<= 11'b10001000101;
		10'd829: y<= 11'b10001000111;
		10'd830: y<= 11'b10001001001;
		10'd831: y<= 11'b10001001100;
		10'd832: y<= 11'b10001001110;
		10'd833: y<= 11'b10001010000;
		10'd834: y<= 11'b10001010011;
		10'd835: y<= 11'b10001010101;
		10'd836: y<= 11'b10001011000;
		10'd837: y<= 11'b10001011010;
		10'd838: y<= 11'b10001011101;
		10'd839: y<= 11'b10001100000;
		10'd840: y<= 11'b10001100010;
		10'd841: y<= 11'b10001100101;
		10'd842: y<= 11'b10001101000;
		10'd843: y<= 11'b10001101011;
		10'd844: y<= 11'b10001101101;
		10'd845: y<= 11'b10001110000;
		10'd846: y<= 11'b10001110011;
		10'd847: y<= 11'b10001110110;
		10'd848: y<= 11'b10001111001;
		10'd849: y<= 11'b10001111100;
		10'd850: y<= 11'b10001111111;
		10'd851: y<= 11'b10010000010;
		10'd852: y<= 11'b10010000101;
		10'd853: y<= 11'b10010001000;
		10'd854: y<= 11'b10010001011;
		10'd855: y<= 11'b10010001110;
		10'd856: y<= 11'b10010010010;
		10'd857: y<= 11'b10010010101;
		10'd858: y<= 11'b10010011000;
		10'd859: y<= 11'b10010011100;
		10'd860: y<= 11'b10010011111;
		10'd861: y<= 11'b10010100010;
		10'd862: y<= 11'b10010100110;
		10'd863: y<= 11'b10010101001;
		10'd864: y<= 11'b10010101101;
		10'd865: y<= 11'b10010110000;
		10'd866: y<= 11'b10010110100;
		10'd867: y<= 11'b10010110111;
		10'd868: y<= 11'b10010111011;
		10'd869: y<= 11'b10010111110;
		10'd870: y<= 11'b10011000010;
		10'd871: y<= 11'b10011000110;
		10'd872: y<= 11'b10011001010;
		10'd873: y<= 11'b10011001101;
		10'd874: y<= 11'b10011010001;
		10'd875: y<= 11'b10011010101;
		10'd876: y<= 11'b10011011001;
		10'd877: y<= 11'b10011011101;
		10'd878: y<= 11'b10011100001;
		10'd879: y<= 11'b10011100100;
		10'd880: y<= 11'b10011101000;
		10'd881: y<= 11'b10011101100;
		10'd882: y<= 11'b10011110000;
		10'd883: y<= 11'b10011110101;
		10'd884: y<= 11'b10011111001;
		10'd885: y<= 11'b10011111101;
		10'd886: y<= 11'b10100000001;
		10'd887: y<= 11'b10100000101;
		10'd888: y<= 11'b10100001001;
		10'd889: y<= 11'b10100001101;
		10'd890: y<= 11'b10100010010;
		10'd891: y<= 11'b10100010110;
		10'd892: y<= 11'b10100011010;
		10'd893: y<= 11'b10100011111;
		10'd894: y<= 11'b10100100011;
		10'd895: y<= 11'b10100100111;
		10'd896: y<= 11'b10100101100;
		10'd897: y<= 11'b10100110000;
		10'd898: y<= 11'b10100110101;
		10'd899: y<= 11'b10100111001;
		10'd900: y<= 11'b10100111110;
		10'd901: y<= 11'b10101000010;
		10'd902: y<= 11'b10101000111;
		10'd903: y<= 11'b10101001100;
		10'd904: y<= 11'b10101010000;
		10'd905: y<= 11'b10101010101;
		10'd906: y<= 11'b10101011010;
		10'd907: y<= 11'b10101011110;
		10'd908: y<= 11'b10101100011;
		10'd909: y<= 11'b10101101000;
		10'd910: y<= 11'b10101101101;
		10'd911: y<= 11'b10101110010;
		10'd912: y<= 11'b10101110110;
		10'd913: y<= 11'b10101111011;
		10'd914: y<= 11'b10110000000;
		10'd915: y<= 11'b10110000101;
		10'd916: y<= 11'b10110001010;
		10'd917: y<= 11'b10110001111;
		10'd918: y<= 11'b10110010100;
		10'd919: y<= 11'b10110011001;
		10'd920: y<= 11'b10110011110;
		10'd921: y<= 11'b10110100011;
		10'd922: y<= 11'b10110101000;
		10'd923: y<= 11'b10110101101;
		10'd924: y<= 11'b10110110010;
		10'd925: y<= 11'b10110111000;
		10'd926: y<= 11'b10110111101;
		10'd927: y<= 11'b10111000010;
		10'd928: y<= 11'b10111000111;
		10'd929: y<= 11'b10111001100;
		10'd930: y<= 11'b10111010010;
		10'd931: y<= 11'b10111010111;
		10'd932: y<= 11'b10111011100;
		10'd933: y<= 11'b10111100001;
		10'd934: y<= 11'b10111100111;
		10'd935: y<= 11'b10111101100;
		10'd936: y<= 11'b10111110010;
		10'd937: y<= 11'b10111110111;
		10'd938: y<= 11'b10111111100;
		10'd939: y<= 11'b11000000010;
		10'd940: y<= 11'b11000000111;
		10'd941: y<= 11'b11000001101;
		10'd942: y<= 11'b11000010010;
		10'd943: y<= 11'b11000011000;
		10'd944: y<= 11'b11000011101;
		10'd945: y<= 11'b11000100011;
		10'd946: y<= 11'b11000101000;
		10'd947: y<= 11'b11000101110;
		10'd948: y<= 11'b11000110100;
		10'd949: y<= 11'b11000111001;
		10'd950: y<= 11'b11000111111;
		10'd951: y<= 11'b11001000101;
		10'd952: y<= 11'b11001001010;
		10'd953: y<= 11'b11001010000;
		10'd954: y<= 11'b11001010110;
		10'd955: y<= 11'b11001011011;
		10'd956: y<= 11'b11001100001;
		10'd957: y<= 11'b11001100111;
		10'd958: y<= 11'b11001101101;
		10'd959: y<= 11'b11001110010;
		10'd960: y<= 11'b11001111000;
		10'd961: y<= 11'b11001111110;
		10'd962: y<= 11'b11010000100;
		10'd963: y<= 11'b11010001010;
		10'd964: y<= 11'b11010001111;
		10'd965: y<= 11'b11010010101;
		10'd966: y<= 11'b11010011011;
		10'd967: y<= 11'b11010100001;
		10'd968: y<= 11'b11010100111;
		10'd969: y<= 11'b11010101101;
		10'd970: y<= 11'b11010110011;
		10'd971: y<= 11'b11010111001;
		10'd972: y<= 11'b11010111111;
		10'd973: y<= 11'b11011000101;
		10'd974: y<= 11'b11011001011;
		10'd975: y<= 11'b11011010001;
		10'd976: y<= 11'b11011010111;
		10'd977: y<= 11'b11011011101;
		10'd978: y<= 11'b11011100011;
		10'd979: y<= 11'b11011101001;
		10'd980: y<= 11'b11011101111;
		10'd981: y<= 11'b11011110101;
		10'd982: y<= 11'b11011111011;
		10'd983: y<= 11'b11100000001;
		10'd984: y<= 11'b11100000111;
		10'd985: y<= 11'b11100001101;
		10'd986: y<= 11'b11100010011;
		10'd987: y<= 11'b11100011010;
		10'd988: y<= 11'b11100100000;
		10'd989: y<= 11'b11100100110;
		10'd990: y<= 11'b11100101100;
		10'd991: y<= 11'b11100110010;
		10'd992: y<= 11'b11100111000;
		10'd993: y<= 11'b11100111110;
		10'd994: y<= 11'b11101000101;
		10'd995: y<= 11'b11101001011;
		10'd996: y<= 11'b11101010001;
		10'd997: y<= 11'b11101010111;
		10'd998: y<= 11'b11101011101;
		10'd999: y<= 11'b11101100100;
		10'd1000: y<= 11'b11101101010;
		10'd1001: y<= 11'b11101110000;
		10'd1002: y<= 11'b11101110110;
		10'd1003: y<= 11'b11101111100;
		10'd1004: y<= 11'b11110000011;
		10'd1005: y<= 11'b11110001001;
		10'd1006: y<= 11'b11110001111;
		10'd1007: y<= 11'b11110010101;
		10'd1008: y<= 11'b11110011100;
		10'd1009: y<= 11'b11110100010;
		10'd1010: y<= 11'b11110101000;
		10'd1011: y<= 11'b11110101110;
		10'd1012: y<= 11'b11110110101;
		10'd1013: y<= 11'b11110111011;
		10'd1014: y<= 11'b11111000001;
		10'd1015: y<= 11'b11111000111;
		10'd1016: y<= 11'b11111001110;
		10'd1017: y<= 11'b11111010100;
		10'd1018: y<= 11'b11111011010;
		10'd1019: y<= 11'b11111100001;
		10'd1020: y<= 11'b11111100111;
		10'd1021: y<= 11'b11111101101;
		10'd1022: y<= 11'b11111110011;
		10'd1023: y<= 11'b11111111010;
     endcase
		//n <= n+1'b1;
	  end
endmodule 