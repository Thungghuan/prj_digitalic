
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:45:04 03/04/2011 
// Design Name: 
// Module Name:    sin_sbox 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module sin_sbox(
input [9:0] sbox_in,
output reg [11:0] sbox_out
);

always @(sbox_in)
	case(sbox_in)		// synopsys full_case parallel_case 
		10'h000: sbox_out= 12'h000;
		10'h001: sbox_out= 12'h006;
		10'h002: sbox_out= 12'h00D;
		10'h003: sbox_out= 12'h013;
		10'h004: sbox_out= 12'h019;
		10'h005: sbox_out= 12'h01F;
		10'h006: sbox_out= 12'h026;
		10'h007: sbox_out= 12'h02C;
		10'h008: sbox_out= 12'h032;
		10'h009: sbox_out= 12'h039;
		10'h00A: sbox_out= 12'h03F;
		10'h00B: sbox_out= 12'h045;
		10'h00C: sbox_out= 12'h04B;
		10'h00D: sbox_out= 12'h052;
		10'h00E: sbox_out= 12'h058;
		10'h00F: sbox_out= 12'h05E;
		10'h010: sbox_out= 12'h064;
		10'h011: sbox_out= 12'h06B;
		10'h012: sbox_out= 12'h071;
		10'h013: sbox_out= 12'h077;
		10'h014: sbox_out= 12'h07D;
		10'h015: sbox_out= 12'h084;
		10'h016: sbox_out= 12'h08A;
		10'h017: sbox_out= 12'h090;
		10'h018: sbox_out= 12'h096;
		10'h019: sbox_out= 12'h09C;
		10'h01A: sbox_out= 12'h0A3;
		10'h01B: sbox_out= 12'h0A9;
		10'h01C: sbox_out= 12'h0AF;
		10'h01D: sbox_out= 12'h0B5;
		10'h01E: sbox_out= 12'h0BB;
		10'h01F: sbox_out= 12'h0C2;
		10'h020: sbox_out= 12'h0C8;
		10'h021: sbox_out= 12'h0CE;
		10'h022: sbox_out= 12'h0D4;
		10'h023: sbox_out= 12'h0DA;
		10'h024: sbox_out= 12'h0E0;
		10'h025: sbox_out= 12'h0E6;
		10'h026: sbox_out= 12'h0ED;
		10'h027: sbox_out= 12'h0F3;
		10'h028: sbox_out= 12'h0F9;
		10'h029: sbox_out= 12'h0FF;
		10'h02A: sbox_out= 12'h105;
		10'h02B: sbox_out= 12'h10B;
		10'h02C: sbox_out= 12'h111;
		10'h02D: sbox_out= 12'h117;
		10'h02E: sbox_out= 12'h11D;
		10'h02F: sbox_out= 12'h123;
		10'h030: sbox_out= 12'h129;
		10'h031: sbox_out= 12'h12F;
		10'h032: sbox_out= 12'h135;
		10'h033: sbox_out= 12'h13B;
		10'h034: sbox_out= 12'h141;
		10'h035: sbox_out= 12'h147;
		10'h036: sbox_out= 12'h14D;
		10'h037: sbox_out= 12'h153;
		10'h038: sbox_out= 12'h159;
		10'h039: sbox_out= 12'h15F;
		10'h03A: sbox_out= 12'h165;
		10'h03B: sbox_out= 12'h16B;
		10'h03C: sbox_out= 12'h171;
		10'h03D: sbox_out= 12'h176;
		10'h03E: sbox_out= 12'h17C;
		10'h03F: sbox_out= 12'h182;
		10'h040: sbox_out= 12'h188;
		10'h041: sbox_out= 12'h18E;
		10'h042: sbox_out= 12'h193;
		10'h043: sbox_out= 12'h199;
		10'h044: sbox_out= 12'h19F;
		10'h045: sbox_out= 12'h1A5;
		10'h046: sbox_out= 12'h1AA;
		10'h047: sbox_out= 12'h1B0;
		10'h048: sbox_out= 12'h1B6;
		10'h049: sbox_out= 12'h1BB;
		10'h04A: sbox_out= 12'h1C1;
		10'h04B: sbox_out= 12'h1C7;
		10'h04C: sbox_out= 12'h1CC;
		10'h04D: sbox_out= 12'h1D2;
		10'h04E: sbox_out= 12'h1D8;
		10'h04F: sbox_out= 12'h1DD;
		10'h050: sbox_out= 12'h1E3;
		10'h051: sbox_out= 12'h1E8;
		10'h052: sbox_out= 12'h1EE;
		10'h053: sbox_out= 12'h1F3;
		10'h054: sbox_out= 12'h1F9;
		10'h055: sbox_out= 12'h1FE;
		10'h056: sbox_out= 12'h204;
		10'h057: sbox_out= 12'h209;
		10'h058: sbox_out= 12'h20E;
		10'h059: sbox_out= 12'h214;
		10'h05A: sbox_out= 12'h219;
		10'h05B: sbox_out= 12'h21F;
		10'h05C: sbox_out= 12'h224;
		10'h05D: sbox_out= 12'h229;
		10'h05E: sbox_out= 12'h22E;
		10'h05F: sbox_out= 12'h234;
		10'h060: sbox_out= 12'h239;
		10'h061: sbox_out= 12'h23E;
		10'h062: sbox_out= 12'h243;
		10'h063: sbox_out= 12'h248;
		10'h064: sbox_out= 12'h24E;
		10'h065: sbox_out= 12'h253;
		10'h066: sbox_out= 12'h258;
		10'h067: sbox_out= 12'h25D;
		10'h068: sbox_out= 12'h262;
		10'h069: sbox_out= 12'h267;
		10'h06A: sbox_out= 12'h26C;
		10'h06B: sbox_out= 12'h271;
		10'h06C: sbox_out= 12'h276;
		10'h06D: sbox_out= 12'h27B;
		10'h06E: sbox_out= 12'h280;
		10'h06F: sbox_out= 12'h285;
		10'h070: sbox_out= 12'h28A;
		10'h071: sbox_out= 12'h28E;
		10'h072: sbox_out= 12'h293;
		10'h073: sbox_out= 12'h298;
		10'h074: sbox_out= 12'h29D;
		10'h075: sbox_out= 12'h2A2;
		10'h076: sbox_out= 12'h2A6;
		10'h077: sbox_out= 12'h2AB;
		10'h078: sbox_out= 12'h2B0;
		10'h079: sbox_out= 12'h2B4;
		10'h07A: sbox_out= 12'h2B9;
		10'h07B: sbox_out= 12'h2BE;
		10'h07C: sbox_out= 12'h2C2;
		10'h07D: sbox_out= 12'h2C7;
		10'h07E: sbox_out= 12'h2CB;
		10'h07F: sbox_out= 12'h2D0;
		10'h080: sbox_out= 12'h2D4;
		10'h081: sbox_out= 12'h2D9;
		10'h082: sbox_out= 12'h2DD;
		10'h083: sbox_out= 12'h2E1;
		10'h084: sbox_out= 12'h2E6;
		10'h085: sbox_out= 12'h2EA;
		10'h086: sbox_out= 12'h2EE;
		10'h087: sbox_out= 12'h2F3;
		10'h088: sbox_out= 12'h2F7;
		10'h089: sbox_out= 12'h2FB;
		10'h08A: sbox_out= 12'h2FF;
		10'h08B: sbox_out= 12'h303;
		10'h08C: sbox_out= 12'h307;
		10'h08D: sbox_out= 12'h30B;
		10'h08E: sbox_out= 12'h310;
		10'h08F: sbox_out= 12'h314;
		10'h090: sbox_out= 12'h318;
		10'h091: sbox_out= 12'h31C;
		10'h092: sbox_out= 12'h31F;
		10'h093: sbox_out= 12'h323;
		10'h094: sbox_out= 12'h327;
		10'h095: sbox_out= 12'h32B;
		10'h096: sbox_out= 12'h32F;
		10'h097: sbox_out= 12'h333;
		10'h098: sbox_out= 12'h336;
		10'h099: sbox_out= 12'h33A;
		10'h09A: sbox_out= 12'h33E;
		10'h09B: sbox_out= 12'h342;
		10'h09C: sbox_out= 12'h345;
		10'h09D: sbox_out= 12'h349;
		10'h09E: sbox_out= 12'h34C;
		10'h09F: sbox_out= 12'h350;
		10'h0A0: sbox_out= 12'h353;
		10'h0A1: sbox_out= 12'h357;
		10'h0A2: sbox_out= 12'h35A;
		10'h0A3: sbox_out= 12'h35E;
		10'h0A4: sbox_out= 12'h361;
		10'h0A5: sbox_out= 12'h364;
		10'h0A6: sbox_out= 12'h368;
		10'h0A7: sbox_out= 12'h36B;
		10'h0A8: sbox_out= 12'h36E;
		10'h0A9: sbox_out= 12'h372;
		10'h0AA: sbox_out= 12'h375;
		10'h0AB: sbox_out= 12'h378;
		10'h0AC: sbox_out= 12'h37B;
		10'h0AD: sbox_out= 12'h37E;
		10'h0AE: sbox_out= 12'h381;
		10'h0AF: sbox_out= 12'h384;
		10'h0B0: sbox_out= 12'h387;
		10'h0B1: sbox_out= 12'h38A;
		10'h0B2: sbox_out= 12'h38D;
		10'h0B3: sbox_out= 12'h390;
		10'h0B4: sbox_out= 12'h393;
		10'h0B5: sbox_out= 12'h395;
		10'h0B6: sbox_out= 12'h398;
		10'h0B7: sbox_out= 12'h39B;
		10'h0B8: sbox_out= 12'h39E;
		10'h0B9: sbox_out= 12'h3A0;
		10'h0BA: sbox_out= 12'h3A3;
		10'h0BB: sbox_out= 12'h3A6;
		10'h0BC: sbox_out= 12'h3A8;
		10'h0BD: sbox_out= 12'h3AB;
		10'h0BE: sbox_out= 12'h3AD;
		10'h0BF: sbox_out= 12'h3B0;
		10'h0C0: sbox_out= 12'h3B2;
		10'h0C1: sbox_out= 12'h3B4;
		10'h0C2: sbox_out= 12'h3B7;
		10'h0C3: sbox_out= 12'h3B9;
		10'h0C4: sbox_out= 12'h3BB;
		10'h0C5: sbox_out= 12'h3BE;
		10'h0C6: sbox_out= 12'h3C0;
		10'h0C7: sbox_out= 12'h3C2;
		10'h0C8: sbox_out= 12'h3C4;
		10'h0C9: sbox_out= 12'h3C6;
		10'h0CA: sbox_out= 12'h3C8;
		10'h0CB: sbox_out= 12'h3CA;
		10'h0CC: sbox_out= 12'h3CC;
		10'h0CD: sbox_out= 12'h3CE;
		10'h0CE: sbox_out= 12'h3D0;
		10'h0CF: sbox_out= 12'h3D2;
		10'h0D0: sbox_out= 12'h3D4;
		10'h0D1: sbox_out= 12'h3D6;
		10'h0D2: sbox_out= 12'h3D7;
		10'h0D3: sbox_out= 12'h3D9;
		10'h0D4: sbox_out= 12'h3DB;
		10'h0D5: sbox_out= 12'h3DD;
		10'h0D6: sbox_out= 12'h3DE;
		10'h0D7: sbox_out= 12'h3E0;
		10'h0D8: sbox_out= 12'h3E1;
		10'h0D9: sbox_out= 12'h3E3;
		10'h0DA: sbox_out= 12'h3E4;
		10'h0DB: sbox_out= 12'h3E6;
		10'h0DC: sbox_out= 12'h3E7;
		10'h0DD: sbox_out= 12'h3E8;
		10'h0DE: sbox_out= 12'h3EA;
		10'h0DF: sbox_out= 12'h3EB;
		10'h0E0: sbox_out= 12'h3EC;
		10'h0E1: sbox_out= 12'h3EE;
		10'h0E2: sbox_out= 12'h3EF;
		10'h0E3: sbox_out= 12'h3F0;
		10'h0E4: sbox_out= 12'h3F1;
		10'h0E5: sbox_out= 12'h3F2;
		10'h0E6: sbox_out= 12'h3F3;
		10'h0E7: sbox_out= 12'h3F4;
		10'h0E8: sbox_out= 12'h3F5;
		10'h0E9: sbox_out= 12'h3F6;
		10'h0EA: sbox_out= 12'h3F7;
		10'h0EB: sbox_out= 12'h3F8;
		10'h0EC: sbox_out= 12'h3F8;
		10'h0ED: sbox_out= 12'h3F9;
		10'h0EE: sbox_out= 12'h3FA;
		10'h0EF: sbox_out= 12'h3FA;
		10'h0F0: sbox_out= 12'h3FB;
		10'h0F1: sbox_out= 12'h3FC;
		10'h0F2: sbox_out= 12'h3FC;
		10'h0F3: sbox_out= 12'h3FD;
		10'h0F4: sbox_out= 12'h3FD;
		10'h0F5: sbox_out= 12'h3FE;
		10'h0F6: sbox_out= 12'h3FE;
		10'h0F7: sbox_out= 12'h3FE;
		10'h0F8: sbox_out= 12'h3FF;
		10'h0F9: sbox_out= 12'h3FF;
		10'h0FA: sbox_out= 12'h3FF;
		10'h0FB: sbox_out= 12'h400;
		10'h0FC: sbox_out= 12'h400;
		10'h0FD: sbox_out= 12'h400;
		10'h0FE: sbox_out= 12'h400;
		10'h0FF: sbox_out= 12'h400;
		10'h100: sbox_out= 12'h400;
		10'h101: sbox_out= 12'h400;
		10'h102: sbox_out= 12'h400;
		10'h103: sbox_out= 12'h400;
		10'h104: sbox_out= 12'h400;
		10'h105: sbox_out= 12'h400;
		10'h106: sbox_out= 12'h3FF;
		10'h107: sbox_out= 12'h3FF;
		10'h108: sbox_out= 12'h3FF;
		10'h109: sbox_out= 12'h3FE;
		10'h10A: sbox_out= 12'h3FE;
		10'h10B: sbox_out= 12'h3FE;
		10'h10C: sbox_out= 12'h3FD;
		10'h10D: sbox_out= 12'h3FD;
		10'h10E: sbox_out= 12'h3FC;
		10'h10F: sbox_out= 12'h3FC;
		10'h110: sbox_out= 12'h3FB;
		10'h111: sbox_out= 12'h3FA;
		10'h112: sbox_out= 12'h3FA;
		10'h113: sbox_out= 12'h3F9;
		10'h114: sbox_out= 12'h3F8;
		10'h115: sbox_out= 12'h3F8;
		10'h116: sbox_out= 12'h3F7;
		10'h117: sbox_out= 12'h3F6;
		10'h118: sbox_out= 12'h3F5;
		10'h119: sbox_out= 12'h3F4;
		10'h11A: sbox_out= 12'h3F3;
		10'h11B: sbox_out= 12'h3F2;
		10'h11C: sbox_out= 12'h3F1;
		10'h11D: sbox_out= 12'h3F0;
		10'h11E: sbox_out= 12'h3EF;
		10'h11F: sbox_out= 12'h3EE;
		10'h120: sbox_out= 12'h3EC;
		10'h121: sbox_out= 12'h3EB;
		10'h122: sbox_out= 12'h3EA;
		10'h123: sbox_out= 12'h3E8;
		10'h124: sbox_out= 12'h3E7;
		10'h125: sbox_out= 12'h3E6;
		10'h126: sbox_out= 12'h3E4;
		10'h127: sbox_out= 12'h3E3;
		10'h128: sbox_out= 12'h3E1;
		10'h129: sbox_out= 12'h3E0;
		10'h12A: sbox_out= 12'h3DE;
		10'h12B: sbox_out= 12'h3DD;
		10'h12C: sbox_out= 12'h3DB;
		10'h12D: sbox_out= 12'h3D9;
		10'h12E: sbox_out= 12'h3D7;
		10'h12F: sbox_out= 12'h3D6;
		10'h130: sbox_out= 12'h3D4;
		10'h131: sbox_out= 12'h3D2;
		10'h132: sbox_out= 12'h3D0;
		10'h133: sbox_out= 12'h3CE;
		10'h134: sbox_out= 12'h3CC;
		10'h135: sbox_out= 12'h3CA;
		10'h136: sbox_out= 12'h3C8;
		10'h137: sbox_out= 12'h3C6;
		10'h138: sbox_out= 12'h3C4;
		10'h139: sbox_out= 12'h3C2;
		10'h13A: sbox_out= 12'h3C0;
		10'h13B: sbox_out= 12'h3BE;
		10'h13C: sbox_out= 12'h3BB;
		10'h13D: sbox_out= 12'h3B9;
		10'h13E: sbox_out= 12'h3B7;
		10'h13F: sbox_out= 12'h3B4;
		10'h140: sbox_out= 12'h3B2;
		10'h141: sbox_out= 12'h3B0;
		10'h142: sbox_out= 12'h3AD;
		10'h143: sbox_out= 12'h3AB;
		10'h144: sbox_out= 12'h3A8;
		10'h145: sbox_out= 12'h3A6;
		10'h146: sbox_out= 12'h3A3;
		10'h147: sbox_out= 12'h3A0;
		10'h148: sbox_out= 12'h39E;
		10'h149: sbox_out= 12'h39B;
		10'h14A: sbox_out= 12'h398;
		10'h14B: sbox_out= 12'h395;
		10'h14C: sbox_out= 12'h393;
		10'h14D: sbox_out= 12'h390;
		10'h14E: sbox_out= 12'h38D;
		10'h14F: sbox_out= 12'h38A;
		10'h150: sbox_out= 12'h387;
		10'h151: sbox_out= 12'h384;
		10'h152: sbox_out= 12'h381;
		10'h153: sbox_out= 12'h37E;
		10'h154: sbox_out= 12'h37B;
		10'h155: sbox_out= 12'h378;
		10'h156: sbox_out= 12'h375;
		10'h157: sbox_out= 12'h372;
		10'h158: sbox_out= 12'h36E;
		10'h159: sbox_out= 12'h36B;
		10'h15A: sbox_out= 12'h368;
		10'h15B: sbox_out= 12'h364;
		10'h15C: sbox_out= 12'h361;
		10'h15D: sbox_out= 12'h35E;
		10'h15E: sbox_out= 12'h35A;
		10'h15F: sbox_out= 12'h357;
		10'h160: sbox_out= 12'h353;
		10'h161: sbox_out= 12'h350;
		10'h162: sbox_out= 12'h34C;
		10'h163: sbox_out= 12'h349;
		10'h164: sbox_out= 12'h345;
		10'h165: sbox_out= 12'h342;
		10'h166: sbox_out= 12'h33E;
		10'h167: sbox_out= 12'h33A;
		10'h168: sbox_out= 12'h336;
		10'h169: sbox_out= 12'h333;
		10'h16A: sbox_out= 12'h32F;
		10'h16B: sbox_out= 12'h32B;
		10'h16C: sbox_out= 12'h327;
		10'h16D: sbox_out= 12'h323;
		10'h16E: sbox_out= 12'h31F;
		10'h16F: sbox_out= 12'h31C;
		10'h170: sbox_out= 12'h318;
		10'h171: sbox_out= 12'h314;
		10'h172: sbox_out= 12'h310;
		10'h173: sbox_out= 12'h30B;
		10'h174: sbox_out= 12'h307;
		10'h175: sbox_out= 12'h303;
		10'h176: sbox_out= 12'h2FF;
		10'h177: sbox_out= 12'h2FB;
		10'h178: sbox_out= 12'h2F7;
		10'h179: sbox_out= 12'h2F3;
		10'h17A: sbox_out= 12'h2EE;
		10'h17B: sbox_out= 12'h2EA;
		10'h17C: sbox_out= 12'h2E6;
		10'h17D: sbox_out= 12'h2E1;
		10'h17E: sbox_out= 12'h2DD;
		10'h17F: sbox_out= 12'h2D9;
		10'h180: sbox_out= 12'h2D4;
		10'h181: sbox_out= 12'h2D0;
		10'h182: sbox_out= 12'h2CB;
		10'h183: sbox_out= 12'h2C7;
		10'h184: sbox_out= 12'h2C2;
		10'h185: sbox_out= 12'h2BE;
		10'h186: sbox_out= 12'h2B9;
		10'h187: sbox_out= 12'h2B4;
		10'h188: sbox_out= 12'h2B0;
		10'h189: sbox_out= 12'h2AB;
		10'h18A: sbox_out= 12'h2A6;
		10'h18B: sbox_out= 12'h2A2;
		10'h18C: sbox_out= 12'h29D;
		10'h18D: sbox_out= 12'h298;
		10'h18E: sbox_out= 12'h293;
		10'h18F: sbox_out= 12'h28E;
		10'h190: sbox_out= 12'h28A;
		10'h191: sbox_out= 12'h285;
		10'h192: sbox_out= 12'h280;
		10'h193: sbox_out= 12'h27B;
		10'h194: sbox_out= 12'h276;
		10'h195: sbox_out= 12'h271;
		10'h196: sbox_out= 12'h26C;
		10'h197: sbox_out= 12'h267;
		10'h198: sbox_out= 12'h262;
		10'h199: sbox_out= 12'h25D;
		10'h19A: sbox_out= 12'h258;
		10'h19B: sbox_out= 12'h253;
		10'h19C: sbox_out= 12'h24E;
		10'h19D: sbox_out= 12'h248;
		10'h19E: sbox_out= 12'h243;
		10'h19F: sbox_out= 12'h23E;
		10'h1A0: sbox_out= 12'h239;
		10'h1A1: sbox_out= 12'h234;
		10'h1A2: sbox_out= 12'h22E;
		10'h1A3: sbox_out= 12'h229;
		10'h1A4: sbox_out= 12'h224;
		10'h1A5: sbox_out= 12'h21F;
		10'h1A6: sbox_out= 12'h219;
		10'h1A7: sbox_out= 12'h214;
		10'h1A8: sbox_out= 12'h20E;
		10'h1A9: sbox_out= 12'h209;
		10'h1AA: sbox_out= 12'h204;
		10'h1AB: sbox_out= 12'h1FE;
		10'h1AC: sbox_out= 12'h1F9;
		10'h1AD: sbox_out= 12'h1F3;
		10'h1AE: sbox_out= 12'h1EE;
		10'h1AF: sbox_out= 12'h1E8;
		10'h1B0: sbox_out= 12'h1E3;
		10'h1B1: sbox_out= 12'h1DD;
		10'h1B2: sbox_out= 12'h1D8;
		10'h1B3: sbox_out= 12'h1D2;
		10'h1B4: sbox_out= 12'h1CC;
		10'h1B5: sbox_out= 12'h1C7;
		10'h1B6: sbox_out= 12'h1C1;
		10'h1B7: sbox_out= 12'h1BB;
		10'h1B8: sbox_out= 12'h1B6;
		10'h1B9: sbox_out= 12'h1B0;
		10'h1BA: sbox_out= 12'h1AA;
		10'h1BB: sbox_out= 12'h1A5;
		10'h1BC: sbox_out= 12'h19F;
		10'h1BD: sbox_out= 12'h199;
		10'h1BE: sbox_out= 12'h193;
		10'h1BF: sbox_out= 12'h18E;
		10'h1C0: sbox_out= 12'h188;
		10'h1C1: sbox_out= 12'h182;
		10'h1C2: sbox_out= 12'h17C;
		10'h1C3: sbox_out= 12'h176;
		10'h1C4: sbox_out= 12'h171;
		10'h1C5: sbox_out= 12'h16B;
		10'h1C6: sbox_out= 12'h165;
		10'h1C7: sbox_out= 12'h15F;
		10'h1C8: sbox_out= 12'h159;
		10'h1C9: sbox_out= 12'h153;
		10'h1CA: sbox_out= 12'h14D;
		10'h1CB: sbox_out= 12'h147;
		10'h1CC: sbox_out= 12'h141;
		10'h1CD: sbox_out= 12'h13B;
		10'h1CE: sbox_out= 12'h135;
		10'h1CF: sbox_out= 12'h12F;
		10'h1D0: sbox_out= 12'h129;
		10'h1D1: sbox_out= 12'h123;
		10'h1D2: sbox_out= 12'h11D;
		10'h1D3: sbox_out= 12'h117;
		10'h1D4: sbox_out= 12'h111;
		10'h1D5: sbox_out= 12'h10B;
		10'h1D6: sbox_out= 12'h105;
		10'h1D7: sbox_out= 12'h0FF;
		10'h1D8: sbox_out= 12'h0F9;
		10'h1D9: sbox_out= 12'h0F3;
		10'h1DA: sbox_out= 12'h0ED;
		10'h1DB: sbox_out= 12'h0E6;
		10'h1DC: sbox_out= 12'h0E0;
		10'h1DD: sbox_out= 12'h0DA;
		10'h1DE: sbox_out= 12'h0D4;
		10'h1DF: sbox_out= 12'h0CE;
		10'h1E0: sbox_out= 12'h0C8;
		10'h1E1: sbox_out= 12'h0C2;
		10'h1E2: sbox_out= 12'h0BB;
		10'h1E3: sbox_out= 12'h0B5;
		10'h1E4: sbox_out= 12'h0AF;
		10'h1E5: sbox_out= 12'h0A9;
		10'h1E6: sbox_out= 12'h0A3;
		10'h1E7: sbox_out= 12'h09C;
		10'h1E8: sbox_out= 12'h096;
		10'h1E9: sbox_out= 12'h090;
		10'h1EA: sbox_out= 12'h08A;
		10'h1EB: sbox_out= 12'h084;
		10'h1EC: sbox_out= 12'h07D;
		10'h1ED: sbox_out= 12'h077;
		10'h1EE: sbox_out= 12'h071;
		10'h1EF: sbox_out= 12'h06B;
		10'h1F0: sbox_out= 12'h064;
		10'h1F1: sbox_out= 12'h05E;
		10'h1F2: sbox_out= 12'h058;
		10'h1F3: sbox_out= 12'h052;
		10'h1F4: sbox_out= 12'h04B;
		10'h1F5: sbox_out= 12'h045;
		10'h1F6: sbox_out= 12'h03F;
		10'h1F7: sbox_out= 12'h039;
		10'h1F8: sbox_out= 12'h032;
		10'h1F9: sbox_out= 12'h02C;
		10'h1FA: sbox_out= 12'h026;
		10'h1FB: sbox_out= 12'h01F;
		10'h1FC: sbox_out= 12'h019;
		10'h1FD: sbox_out= 12'h013;
		10'h1FE: sbox_out= 12'h00D;
		10'h1FF: sbox_out= 12'h006;
		10'h200: sbox_out= 12'h000;
		10'h201: sbox_out= 12'hFFA;
		10'h202: sbox_out= 12'hFF3;
		10'h203: sbox_out= 12'hFED;
		10'h204: sbox_out= 12'hFE7;
		10'h205: sbox_out= 12'hFE1;
		10'h206: sbox_out= 12'hFDA;
		10'h207: sbox_out= 12'hFD4;
		10'h208: sbox_out= 12'hFCE;
		10'h209: sbox_out= 12'hFC7;
		10'h20A: sbox_out= 12'hFC1;
		10'h20B: sbox_out= 12'hFBB;
		10'h20C: sbox_out= 12'hFB5;
		10'h20D: sbox_out= 12'hFAE;
		10'h20E: sbox_out= 12'hFA8;
		10'h20F: sbox_out= 12'hFA2;
		10'h210: sbox_out= 12'hF9C;
		10'h211: sbox_out= 12'hF95;
		10'h212: sbox_out= 12'hF8F;
		10'h213: sbox_out= 12'hF89;
		10'h214: sbox_out= 12'hF83;
		10'h215: sbox_out= 12'hF7C;
		10'h216: sbox_out= 12'hF76;
		10'h217: sbox_out= 12'hF70;
		10'h218: sbox_out= 12'hF6A;
		10'h219: sbox_out= 12'hF64;
		10'h21A: sbox_out= 12'hF5D;
		10'h21B: sbox_out= 12'hF57;
		10'h21C: sbox_out= 12'hF51;
		10'h21D: sbox_out= 12'hF4B;
		10'h21E: sbox_out= 12'hF45;
		10'h21F: sbox_out= 12'hF3E;
		10'h220: sbox_out= 12'hF38;
		10'h221: sbox_out= 12'hF32;
		10'h222: sbox_out= 12'hF2C;
		10'h223: sbox_out= 12'hF26;
		10'h224: sbox_out= 12'hF20;
		10'h225: sbox_out= 12'hF1A;
		10'h226: sbox_out= 12'hF13;
		10'h227: sbox_out= 12'hF0D;
		10'h228: sbox_out= 12'hF07;
		10'h229: sbox_out= 12'hF01;
		10'h22A: sbox_out= 12'hEFB;
		10'h22B: sbox_out= 12'hEF5;
		10'h22C: sbox_out= 12'hEEF;
		10'h22D: sbox_out= 12'hEE9;
		10'h22E: sbox_out= 12'hEE3;
		10'h22F: sbox_out= 12'hEDD;
		10'h230: sbox_out= 12'hED7;
		10'h231: sbox_out= 12'hED1;
		10'h232: sbox_out= 12'hECB;
		10'h233: sbox_out= 12'hEC5;
		10'h234: sbox_out= 12'hEBF;
		10'h235: sbox_out= 12'hEB9;
		10'h236: sbox_out= 12'hEB3;
		10'h237: sbox_out= 12'hEAD;
		10'h238: sbox_out= 12'hEA7;
		10'h239: sbox_out= 12'hEA1;
		10'h23A: sbox_out= 12'hE9B;
		10'h23B: sbox_out= 12'hE95;
		10'h23C: sbox_out= 12'hE8F;
		10'h23D: sbox_out= 12'hE8A;
		10'h23E: sbox_out= 12'hE84;
		10'h23F: sbox_out= 12'hE7E;
		10'h240: sbox_out= 12'hE78;
		10'h241: sbox_out= 12'hE72;
		10'h242: sbox_out= 12'hE6D;
		10'h243: sbox_out= 12'hE67;
		10'h244: sbox_out= 12'hE61;
		10'h245: sbox_out= 12'hE5B;
		10'h246: sbox_out= 12'hE56;
		10'h247: sbox_out= 12'hE50;
		10'h248: sbox_out= 12'hE4A;
		10'h249: sbox_out= 12'hE45;
		10'h24A: sbox_out= 12'hE3F;
		10'h24B: sbox_out= 12'hE39;
		10'h24C: sbox_out= 12'hE34;
		10'h24D: sbox_out= 12'hE2E;
		10'h24E: sbox_out= 12'hE28;
		10'h24F: sbox_out= 12'hE23;
		10'h250: sbox_out= 12'hE1D;
		10'h251: sbox_out= 12'hE18;
		10'h252: sbox_out= 12'hE12;
		10'h253: sbox_out= 12'hE0D;
		10'h254: sbox_out= 12'hE07;
		10'h255: sbox_out= 12'hE02;
		10'h256: sbox_out= 12'hDFC;
		10'h257: sbox_out= 12'hDF7;
		10'h258: sbox_out= 12'hDF2;
		10'h259: sbox_out= 12'hDEC;
		10'h25A: sbox_out= 12'hDE7;
		10'h25B: sbox_out= 12'hDE1;
		10'h25C: sbox_out= 12'hDDC;
		10'h25D: sbox_out= 12'hDD7;
		10'h25E: sbox_out= 12'hDD2;
		10'h25F: sbox_out= 12'hDCC;
		10'h260: sbox_out= 12'hDC7;
		10'h261: sbox_out= 12'hDC2;
		10'h262: sbox_out= 12'hDBD;
		10'h263: sbox_out= 12'hDB8;
		10'h264: sbox_out= 12'hDB2;
		10'h265: sbox_out= 12'hDAD;
		10'h266: sbox_out= 12'hDA8;
		10'h267: sbox_out= 12'hDA3;
		10'h268: sbox_out= 12'hD9E;
		10'h269: sbox_out= 12'hD99;
		10'h26A: sbox_out= 12'hD94;
		10'h26B: sbox_out= 12'hD8F;
		10'h26C: sbox_out= 12'hD8A;
		10'h26D: sbox_out= 12'hD85;
		10'h26E: sbox_out= 12'hD80;
		10'h26F: sbox_out= 12'hD7B;
		10'h270: sbox_out= 12'hD76;
		10'h271: sbox_out= 12'hD72;
		10'h272: sbox_out= 12'hD6D;
		10'h273: sbox_out= 12'hD68;
		10'h274: sbox_out= 12'hD63;
		10'h275: sbox_out= 12'hD5E;
		10'h276: sbox_out= 12'hD5A;
		10'h277: sbox_out= 12'hD55;
		10'h278: sbox_out= 12'hD50;
		10'h279: sbox_out= 12'hD4C;
		10'h27A: sbox_out= 12'hD47;
		10'h27B: sbox_out= 12'hD42;
		10'h27C: sbox_out= 12'hD3E;
		10'h27D: sbox_out= 12'hD39;
		10'h27E: sbox_out= 12'hD35;
		10'h27F: sbox_out= 12'hD30;
		10'h280: sbox_out= 12'hD2C;
		10'h281: sbox_out= 12'hD27;
		10'h282: sbox_out= 12'hD23;
		10'h283: sbox_out= 12'hD1F;
		10'h284: sbox_out= 12'hD1A;
		10'h285: sbox_out= 12'hD16;
		10'h286: sbox_out= 12'hD12;
		10'h287: sbox_out= 12'hD0D;
		10'h288: sbox_out= 12'hD09;
		10'h289: sbox_out= 12'hD05;
		10'h28A: sbox_out= 12'hD01;
		10'h28B: sbox_out= 12'hCFD;
		10'h28C: sbox_out= 12'hCF9;
		10'h28D: sbox_out= 12'hCF5;
		10'h28E: sbox_out= 12'hCF0;
		10'h28F: sbox_out= 12'hCEC;
		10'h290: sbox_out= 12'hCE8;
		10'h291: sbox_out= 12'hCE4;
		10'h292: sbox_out= 12'hCE1;
		10'h293: sbox_out= 12'hCDD;
		10'h294: sbox_out= 12'hCD9;
		10'h295: sbox_out= 12'hCD5;
		10'h296: sbox_out= 12'hCD1;
		10'h297: sbox_out= 12'hCCD;
		10'h298: sbox_out= 12'hCCA;
		10'h299: sbox_out= 12'hCC6;
		10'h29A: sbox_out= 12'hCC2;
		10'h29B: sbox_out= 12'hCBE;
		10'h29C: sbox_out= 12'hCBB;
		10'h29D: sbox_out= 12'hCB7;
		10'h29E: sbox_out= 12'hCB4;
		10'h29F: sbox_out= 12'hCB0;
		10'h2A0: sbox_out= 12'hCAD;
		10'h2A1: sbox_out= 12'hCA9;
		10'h2A2: sbox_out= 12'hCA6;
		10'h2A3: sbox_out= 12'hCA2;
		10'h2A4: sbox_out= 12'hC9F;
		10'h2A5: sbox_out= 12'hC9C;
		10'h2A6: sbox_out= 12'hC98;
		10'h2A7: sbox_out= 12'hC95;
		10'h2A8: sbox_out= 12'hC92;
		10'h2A9: sbox_out= 12'hC8E;
		10'h2AA: sbox_out= 12'hC8B;
		10'h2AB: sbox_out= 12'hC88;
		10'h2AC: sbox_out= 12'hC85;
		10'h2AD: sbox_out= 12'hC82;
		10'h2AE: sbox_out= 12'hC7F;
		10'h2AF: sbox_out= 12'hC7C;
		10'h2B0: sbox_out= 12'hC79;
		10'h2B1: sbox_out= 12'hC76;
		10'h2B2: sbox_out= 12'hC73;
		10'h2B3: sbox_out= 12'hC70;
		10'h2B4: sbox_out= 12'hC6D;
		10'h2B5: sbox_out= 12'hC6B;
		10'h2B6: sbox_out= 12'hC68;
		10'h2B7: sbox_out= 12'hC65;
		10'h2B8: sbox_out= 12'hC62;
		10'h2B9: sbox_out= 12'hC60;
		10'h2BA: sbox_out= 12'hC5D;
		10'h2BB: sbox_out= 12'hC5A;
		10'h2BC: sbox_out= 12'hC58;
		10'h2BD: sbox_out= 12'hC55;
		10'h2BE: sbox_out= 12'hC53;
		10'h2BF: sbox_out= 12'hC50;
		10'h2C0: sbox_out= 12'hC4E;
		10'h2C1: sbox_out= 12'hC4C;
		10'h2C2: sbox_out= 12'hC49;
		10'h2C3: sbox_out= 12'hC47;
		10'h2C4: sbox_out= 12'hC45;
		10'h2C5: sbox_out= 12'hC42;
		10'h2C6: sbox_out= 12'hC40;
		10'h2C7: sbox_out= 12'hC3E;
		10'h2C8: sbox_out= 12'hC3C;
		10'h2C9: sbox_out= 12'hC3A;
		10'h2CA: sbox_out= 12'hC38;
		10'h2CB: sbox_out= 12'hC36;
		10'h2CC: sbox_out= 12'hC34;
		10'h2CD: sbox_out= 12'hC32;
		10'h2CE: sbox_out= 12'hC30;
		10'h2CF: sbox_out= 12'hC2E;
		10'h2D0: sbox_out= 12'hC2C;
		10'h2D1: sbox_out= 12'hC2A;
		10'h2D2: sbox_out= 12'hC29;
		10'h2D3: sbox_out= 12'hC27;
		10'h2D4: sbox_out= 12'hC25;
		10'h2D5: sbox_out= 12'hC23;
		10'h2D6: sbox_out= 12'hC22;
		10'h2D7: sbox_out= 12'hC20;
		10'h2D8: sbox_out= 12'hC1F;
		10'h2D9: sbox_out= 12'hC1D;
		10'h2DA: sbox_out= 12'hC1C;
		10'h2DB: sbox_out= 12'hC1A;
		10'h2DC: sbox_out= 12'hC19;
		10'h2DD: sbox_out= 12'hC18;
		10'h2DE: sbox_out= 12'hC16;
		10'h2DF: sbox_out= 12'hC15;
		10'h2E0: sbox_out= 12'hC14;
		10'h2E1: sbox_out= 12'hC12;
		10'h2E2: sbox_out= 12'hC11;
		10'h2E3: sbox_out= 12'hC10;
		10'h2E4: sbox_out= 12'hC0F;
		10'h2E5: sbox_out= 12'hC0E;
		10'h2E6: sbox_out= 12'hC0D;
		10'h2E7: sbox_out= 12'hC0C;
		10'h2E8: sbox_out= 12'hC0B;
		10'h2E9: sbox_out= 12'hC0A;
		10'h2EA: sbox_out= 12'hC09;
		10'h2EB: sbox_out= 12'hC08;
		10'h2EC: sbox_out= 12'hC08;
		10'h2ED: sbox_out= 12'hC07;
		10'h2EE: sbox_out= 12'hC06;
		10'h2EF: sbox_out= 12'hC06;
		10'h2F0: sbox_out= 12'hC05;
		10'h2F1: sbox_out= 12'hC04;
		10'h2F2: sbox_out= 12'hC04;
		10'h2F3: sbox_out= 12'hC03;
		10'h2F4: sbox_out= 12'hC03;
		10'h2F5: sbox_out= 12'hC02;
		10'h2F6: sbox_out= 12'hC02;
		10'h2F7: sbox_out= 12'hC02;
		10'h2F8: sbox_out= 12'hC01;
		10'h2F9: sbox_out= 12'hC01;
		10'h2FA: sbox_out= 12'hC01;
		10'h2FB: sbox_out= 12'hC00;
		10'h2FC: sbox_out= 12'hC00;
		10'h2FD: sbox_out= 12'hC00;
		10'h2FE: sbox_out= 12'hC00;
		10'h2FF: sbox_out= 12'hC00;
		10'h300: sbox_out= 12'hC00;
		10'h301: sbox_out= 12'hC00;
		10'h302: sbox_out= 12'hC00;
		10'h303: sbox_out= 12'hC00;
		10'h304: sbox_out= 12'hC00;
		10'h305: sbox_out= 12'hC00;
		10'h306: sbox_out= 12'hC01;
		10'h307: sbox_out= 12'hC01;
		10'h308: sbox_out= 12'hC01;
		10'h309: sbox_out= 12'hC02;
		10'h30A: sbox_out= 12'hC02;
		10'h30B: sbox_out= 12'hC02;
		10'h30C: sbox_out= 12'hC03;
		10'h30D: sbox_out= 12'hC03;
		10'h30E: sbox_out= 12'hC04;
		10'h30F: sbox_out= 12'hC04;
		10'h310: sbox_out= 12'hC05;
		10'h311: sbox_out= 12'hC06;
		10'h312: sbox_out= 12'hC06;
		10'h313: sbox_out= 12'hC07;
		10'h314: sbox_out= 12'hC08;
		10'h315: sbox_out= 12'hC08;
		10'h316: sbox_out= 12'hC09;
		10'h317: sbox_out= 12'hC0A;
		10'h318: sbox_out= 12'hC0B;
		10'h319: sbox_out= 12'hC0C;
		10'h31A: sbox_out= 12'hC0D;
		10'h31B: sbox_out= 12'hC0E;
		10'h31C: sbox_out= 12'hC0F;
		10'h31D: sbox_out= 12'hC10;
		10'h31E: sbox_out= 12'hC11;
		10'h31F: sbox_out= 12'hC12;
		10'h320: sbox_out= 12'hC14;
		10'h321: sbox_out= 12'hC15;
		10'h322: sbox_out= 12'hC16;
		10'h323: sbox_out= 12'hC18;
		10'h324: sbox_out= 12'hC19;
		10'h325: sbox_out= 12'hC1A;
		10'h326: sbox_out= 12'hC1C;
		10'h327: sbox_out= 12'hC1D;
		10'h328: sbox_out= 12'hC1F;
		10'h329: sbox_out= 12'hC20;
		10'h32A: sbox_out= 12'hC22;
		10'h32B: sbox_out= 12'hC23;
		10'h32C: sbox_out= 12'hC25;
		10'h32D: sbox_out= 12'hC27;
		10'h32E: sbox_out= 12'hC29;
		10'h32F: sbox_out= 12'hC2A;
		10'h330: sbox_out= 12'hC2C;
		10'h331: sbox_out= 12'hC2E;
		10'h332: sbox_out= 12'hC30;
		10'h333: sbox_out= 12'hC32;
		10'h334: sbox_out= 12'hC34;
		10'h335: sbox_out= 12'hC36;
		10'h336: sbox_out= 12'hC38;
		10'h337: sbox_out= 12'hC3A;
		10'h338: sbox_out= 12'hC3C;
		10'h339: sbox_out= 12'hC3E;
		10'h33A: sbox_out= 12'hC40;
		10'h33B: sbox_out= 12'hC42;
		10'h33C: sbox_out= 12'hC45;
		10'h33D: sbox_out= 12'hC47;
		10'h33E: sbox_out= 12'hC49;
		10'h33F: sbox_out= 12'hC4C;
		10'h340: sbox_out= 12'hC4E;
		10'h341: sbox_out= 12'hC50;
		10'h342: sbox_out= 12'hC53;
		10'h343: sbox_out= 12'hC55;
		10'h344: sbox_out= 12'hC58;
		10'h345: sbox_out= 12'hC5A;
		10'h346: sbox_out= 12'hC5D;
		10'h347: sbox_out= 12'hC60;
		10'h348: sbox_out= 12'hC62;
		10'h349: sbox_out= 12'hC65;
		10'h34A: sbox_out= 12'hC68;
		10'h34B: sbox_out= 12'hC6B;
		10'h34C: sbox_out= 12'hC6D;
		10'h34D: sbox_out= 12'hC70;
		10'h34E: sbox_out= 12'hC73;
		10'h34F: sbox_out= 12'hC76;
		10'h350: sbox_out= 12'hC79;
		10'h351: sbox_out= 12'hC7C;
		10'h352: sbox_out= 12'hC7F;
		10'h353: sbox_out= 12'hC82;
		10'h354: sbox_out= 12'hC85;
		10'h355: sbox_out= 12'hC88;
		10'h356: sbox_out= 12'hC8B;
		10'h357: sbox_out= 12'hC8E;
		10'h358: sbox_out= 12'hC92;
		10'h359: sbox_out= 12'hC95;
		10'h35A: sbox_out= 12'hC98;
		10'h35B: sbox_out= 12'hC9C;
		10'h35C: sbox_out= 12'hC9F;
		10'h35D: sbox_out= 12'hCA2;
		10'h35E: sbox_out= 12'hCA6;
		10'h35F: sbox_out= 12'hCA9;
		10'h360: sbox_out= 12'hCAD;
		10'h361: sbox_out= 12'hCB0;
		10'h362: sbox_out= 12'hCB4;
		10'h363: sbox_out= 12'hCB7;
		10'h364: sbox_out= 12'hCBB;
		10'h365: sbox_out= 12'hCBE;
		10'h366: sbox_out= 12'hCC2;
		10'h367: sbox_out= 12'hCC6;
		10'h368: sbox_out= 12'hCCA;
		10'h369: sbox_out= 12'hCCD;
		10'h36A: sbox_out= 12'hCD1;
		10'h36B: sbox_out= 12'hCD5;
		10'h36C: sbox_out= 12'hCD9;
		10'h36D: sbox_out= 12'hCDD;
		10'h36E: sbox_out= 12'hCE1;
		10'h36F: sbox_out= 12'hCE4;
		10'h370: sbox_out= 12'hCE8;
		10'h371: sbox_out= 12'hCEC;
		10'h372: sbox_out= 12'hCF0;
		10'h373: sbox_out= 12'hCF5;
		10'h374: sbox_out= 12'hCF9;
		10'h375: sbox_out= 12'hCFD;
		10'h376: sbox_out= 12'hD01;
		10'h377: sbox_out= 12'hD05;
		10'h378: sbox_out= 12'hD09;
		10'h379: sbox_out= 12'hD0D;
		10'h37A: sbox_out= 12'hD12;
		10'h37B: sbox_out= 12'hD16;
		10'h37C: sbox_out= 12'hD1A;
		10'h37D: sbox_out= 12'hD1F;
		10'h37E: sbox_out= 12'hD23;
		10'h37F: sbox_out= 12'hD27;
		10'h380: sbox_out= 12'hD2C;
		10'h381: sbox_out= 12'hD30;
		10'h382: sbox_out= 12'hD35;
		10'h383: sbox_out= 12'hD39;
		10'h384: sbox_out= 12'hD3E;
		10'h385: sbox_out= 12'hD42;
		10'h386: sbox_out= 12'hD47;
		10'h387: sbox_out= 12'hD4C;
		10'h388: sbox_out= 12'hD50;
		10'h389: sbox_out= 12'hD55;
		10'h38A: sbox_out= 12'hD5A;
		10'h38B: sbox_out= 12'hD5E;
		10'h38C: sbox_out= 12'hD63;
		10'h38D: sbox_out= 12'hD68;
		10'h38E: sbox_out= 12'hD6D;
		10'h38F: sbox_out= 12'hD72;
		10'h390: sbox_out= 12'hD76;
		10'h391: sbox_out= 12'hD7B;
		10'h392: sbox_out= 12'hD80;
		10'h393: sbox_out= 12'hD85;
		10'h394: sbox_out= 12'hD8A;
		10'h395: sbox_out= 12'hD8F;
		10'h396: sbox_out= 12'hD94;
		10'h397: sbox_out= 12'hD99;
		10'h398: sbox_out= 12'hD9E;
		10'h399: sbox_out= 12'hDA3;
		10'h39A: sbox_out= 12'hDA8;
		10'h39B: sbox_out= 12'hDAD;
		10'h39C: sbox_out= 12'hDB2;
		10'h39D: sbox_out= 12'hDB8;
		10'h39E: sbox_out= 12'hDBD;
		10'h39F: sbox_out= 12'hDC2;
		10'h3A0: sbox_out= 12'hDC7;
		10'h3A1: sbox_out= 12'hDCC;
		10'h3A2: sbox_out= 12'hDD2;
		10'h3A3: sbox_out= 12'hDD7;
		10'h3A4: sbox_out= 12'hDDC;
		10'h3A5: sbox_out= 12'hDE1;
		10'h3A6: sbox_out= 12'hDE7;
		10'h3A7: sbox_out= 12'hDEC;
		10'h3A8: sbox_out= 12'hDF2;
		10'h3A9: sbox_out= 12'hDF7;
		10'h3AA: sbox_out= 12'hDFC;
		10'h3AB: sbox_out= 12'hE02;
		10'h3AC: sbox_out= 12'hE07;
		10'h3AD: sbox_out= 12'hE0D;
		10'h3AE: sbox_out= 12'hE12;
		10'h3AF: sbox_out= 12'hE18;
		10'h3B0: sbox_out= 12'hE1D;
		10'h3B1: sbox_out= 12'hE23;
		10'h3B2: sbox_out= 12'hE28;
		10'h3B3: sbox_out= 12'hE2E;
		10'h3B4: sbox_out= 12'hE34;
		10'h3B5: sbox_out= 12'hE39;
		10'h3B6: sbox_out= 12'hE3F;
		10'h3B7: sbox_out= 12'hE45;
		10'h3B8: sbox_out= 12'hE4A;
		10'h3B9: sbox_out= 12'hE50;
		10'h3BA: sbox_out= 12'hE56;
		10'h3BB: sbox_out= 12'hE5B;
		10'h3BC: sbox_out= 12'hE61;
		10'h3BD: sbox_out= 12'hE67;
		10'h3BE: sbox_out= 12'hE6D;
		10'h3BF: sbox_out= 12'hE72;
		10'h3C0: sbox_out= 12'hE78;
		10'h3C1: sbox_out= 12'hE7E;
		10'h3C2: sbox_out= 12'hE84;
		10'h3C3: sbox_out= 12'hE8A;
		10'h3C4: sbox_out= 12'hE8F;
		10'h3C5: sbox_out= 12'hE95;
		10'h3C6: sbox_out= 12'hE9B;
		10'h3C7: sbox_out= 12'hEA1;
		10'h3C8: sbox_out= 12'hEA7;
		10'h3C9: sbox_out= 12'hEAD;
		10'h3CA: sbox_out= 12'hEB3;
		10'h3CB: sbox_out= 12'hEB9;
		10'h3CC: sbox_out= 12'hEBF;
		10'h3CD: sbox_out= 12'hEC5;
		10'h3CE: sbox_out= 12'hECB;
		10'h3CF: sbox_out= 12'hED1;
		10'h3D0: sbox_out= 12'hED7;
		10'h3D1: sbox_out= 12'hEDD;
		10'h3D2: sbox_out= 12'hEE3;
		10'h3D3: sbox_out= 12'hEE9;
		10'h3D4: sbox_out= 12'hEEF;
		10'h3D5: sbox_out= 12'hEF5;
		10'h3D6: sbox_out= 12'hEFB;
		10'h3D7: sbox_out= 12'hF01;
		10'h3D8: sbox_out= 12'hF07;
		10'h3D9: sbox_out= 12'hF0D;
		10'h3DA: sbox_out= 12'hF13;
		10'h3DB: sbox_out= 12'hF1A;
		10'h3DC: sbox_out= 12'hF20;
		10'h3DD: sbox_out= 12'hF26;
		10'h3DE: sbox_out= 12'hF2C;
		10'h3DF: sbox_out= 12'hF32;
		10'h3E0: sbox_out= 12'hF38;
		10'h3E1: sbox_out= 12'hF3E;
		10'h3E2: sbox_out= 12'hF45;
		10'h3E3: sbox_out= 12'hF4B;
		10'h3E4: sbox_out= 12'hF51;
		10'h3E5: sbox_out= 12'hF57;
		10'h3E6: sbox_out= 12'hF5D;
		10'h3E7: sbox_out= 12'hF64;
		10'h3E8: sbox_out= 12'hF6A;
		10'h3E9: sbox_out= 12'hF70;
		10'h3EA: sbox_out= 12'hF76;
		10'h3EB: sbox_out= 12'hF7C;
		10'h3EC: sbox_out= 12'hF83;
		10'h3ED: sbox_out= 12'hF89;
		10'h3EE: sbox_out= 12'hF8F;
		10'h3EF: sbox_out= 12'hF95;
		10'h3F0: sbox_out= 12'hF9C;
		10'h3F1: sbox_out= 12'hFA2;
		10'h3F2: sbox_out= 12'hFA8;
		10'h3F3: sbox_out= 12'hFAE;
		10'h3F4: sbox_out= 12'hFB5;
		10'h3F5: sbox_out= 12'hFBB;
		10'h3F6: sbox_out= 12'hFC1;
		10'h3F7: sbox_out= 12'hFC7;
		10'h3F8: sbox_out= 12'hFCE;
		10'h3F9: sbox_out= 12'hFD4;
		10'h3FA: sbox_out= 12'hFDA;
		10'h3FB: sbox_out= 12'hFE1;
		10'h3FC: sbox_out= 12'hFE7;
		10'h3FD: sbox_out= 12'hFED;
		10'h3FE: sbox_out= 12'hFF3;
		10'h3FF: sbox_out= 12'hFFA;

	endcase

endmodule
